--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
--	Grupo de Apoio ao Projeto de Hardware  - GAPH
--	Projeto X10GiGA - FINEP/PUCRS/TERACOM
--
--	M�dulo:	Mem�ria - Gerador de Frames - Prototipa��o
--	Autor:	Jeferson Camargo de Oliveira
--
-- 	FRAME:	0003
-- 	RAMB:	03
-- 	CONJ:	A
--
--	M�dulo gerado em 17 de July de 2008 �s 16h55min pelo
--	programa gerador de frames OTN do projeto X10GiGA.
--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

----Pragma translate_off
library unisim ;
use unisim.vcomponents.all ;
----Pragma translate_on

entity FRAME0003_A3 is
port(
		addr	: in  std_logic_vector(9 downto 0);	-- Barramento de endere�os da porta
		clk		: in  std_logic;					-- Entrada de clock para a porta
		dout	: out std_logic_vector(15 downto 0)	-- Sa�da de dados da porta
	);
end FRAME0003_A3;

architecture FRAME0003_A3 of FRAME0003_A3 is

	signal addrin	: std_logic_vector(9 downto 0);
	signal clkin	: std_logic;
	signal doutout	: std_logic_vector(15 downto 0);

	component RAMB16_S18 is
	generic(
		WRITE_MODE : string;
		INIT_00,INIT_01,INIT_02,INIT_03,INIT_04,INIT_05,INIT_06,INIT_07,
		INIT_08,INIT_09,INIT_0A,INIT_0B,INIT_0C,INIT_0D,INIT_0E,INIT_0F,
		INIT_10,INIT_11,INIT_12,INIT_13,INIT_14,INIT_15,INIT_16,INIT_17,
		INIT_18,INIT_19,INIT_1A,INIT_1B,INIT_1C,INIT_1D,INIT_1E,INIT_1F,
		INIT_20,INIT_21,INIT_22,INIT_23,INIT_24,INIT_25,INIT_26,INIT_27,
		INIT_28,INIT_29,INIT_2A,INIT_2B,INIT_2C,INIT_2D,INIT_2E,INIT_2F,
		INIT_30,INIT_31,INIT_32,INIT_33,INIT_34,INIT_35,INIT_36,INIT_37,
		INIT_38,INIT_39,INIT_3A,INIT_3B,INIT_3C,INIT_3D,INIT_3E,INIT_3F : bit_vector
	);
	port(
		DO   : out std_logic_vector(15 downto 0);	-- Port 16-bit Data Output
		DOP  : out std_logic_vector(1  downto 0);	-- Port 2-bit Parity Output
		ADDR : in  std_logic_vector(9  downto 0); 	-- Port 10-bit Address Input
		CLK  : in  std_logic;			 			-- Port Clock
		DI   : in  std_logic_vector(15 downto 0); 	-- Port 16-bit Data Input
		DIP  : in  std_logic_vector(1  downto 0); 	-- Port 2-bit parity Input
		EN   : in  std_logic;			 			-- Port RAM Enable Input
		SSR  : in  std_logic;			 			-- Port Synchronous Set/Reset Input
		WE   : in  std_logic			 			-- Port Write Enable Input
	);
	end component;

begin

	addrin <= addr;
	clkin  <= clk;
	dout   <= doutout;

	-- FRAME0003_RAMB03 instantiation
	FRAME0003_RAMB03 : RAMB16_S18
	generic map (

		-- The following generics are only necessary if you wish to change the default behavior.
		WRITE_MODE => "NO_CHANGE", 	-- WRITE_FIRST, READ_FIRST or NO_CHANGE

		-- The following generic INIT_xx declarations are only necessary
		-- if you wish to change the initial contents of the RAM to anything
		-- other than all zero's.
		INIT_00 => x"99C3B0AB2F0D91F6F250F2115EC8E33099B7D02ACCE8FAA87EE73A3477E7FCFF",
		INIT_01 => x"D5E5D4D70D7634D785A1ADE9033418712C3B889CEF925D92AF2B2A19AAC6B145",
		INIT_02 => x"1BDB703E531E3D36FA18BE2263810574D3A4B4F07D8CC3EF89A4ECEA3ECC49C8",
		INIT_03 => x"00841B9318961FC358928B0413C781972FE8379CA063A12D2E8AD19ECBD48197",
		INIT_04 => x"020E459BF8F7E69FEDA9E08EDF13BF69E6E82C841D6CE4846BA7FB7E7710D129",
		INIT_05 => x"34674A9783007AB1C4364435F21555A8B6F2E3EA5824CF48A032E219C2152F07",
		INIT_06 => x"001F66D21D4B6AE652E43DF1E7F6814E6C9B7A48323069E5B924FCBD5C26BEE4",
		INIT_07 => x"B4752A8081A89603EB5C95CA383863D5463ED676AFBB6A2B0DE824612BD5F186",
		INIT_08 => x"231E1314644BF78A2CF1C02D3B876C06556A785ACEB77DE2D9AD3E61C3D3BFC9",
		INIT_09 => x"171CD1B6DBCC7CAF034A7EE91C5A8920995951A44314EFE8C740B4D17544E348",
		INIT_0A => x"0B0F5EFFAD5483E2782E45518161D4B1BD511D784039112D2ED24CD3FDE0A0A0",
		INIT_0B => x"5C175802513A0E348C6652206C7C47E695F7BE216E2F988A94CB440508BD2E48",
		INIT_0C => x"429A166C87B2B339510B1C910454B9BE5779A3B71C186E92519536BDE4879323",
		INIT_0D => x"3C843257D989DD65B4FD0D40B329FF9C3F7A13607C423A14DA2B5CCF20D921AC",
		INIT_0E => x"AD3FEC7635D92F52323704923525B78595A74FA8224A5A5EE86E4A5BB0E170C1",
		INIT_0F => x"BC837C4468B72A3E002C4F68F54A42B5EA0830D32875006E466DC367AA78681E",
		INIT_10 => x"E97C3F955C3B215019F011428F68875550A5B10F7AA061CE5FE7B13C79ADAF9B",
		INIT_11 => x"84E138D7C01DFC1625716219897CD4643F600D8A64AE558C8362B18FAE6BE199",
		INIT_12 => x"318DE7F751423A418D680B0CA849E468BE3B08590AFD2CC99D7004C3CF7570BA",
		INIT_13 => x"13BB9B062DF1A91863450FB24EB53DC05711B4282C1F32A1D82EFC122BBD608B",
		INIT_14 => x"938AA734D5F1129E57E271D7BFC317E685A4638BC46F50032D440F87DE4B8612",
		INIT_15 => x"0F74C42D40E3816669B9A864E57D62858E726D075C04CBD1C3DB2C338A55C19B",
		INIT_16 => x"BFC0C802C6760EAEBBF5592D3E0ED02E404F88669706A808FFB97A3806C44A7A",
		INIT_17 => x"0840433424B0FC37A74624183AC4F60E0B4E01D2032BCA60EAFCF682F36FE4B4",
		INIT_18 => x"8E462F396A8055ABA4F2137E0B9360A5C06A1F1D886AB4886EA81E67511992B2",
		INIT_19 => x"F1C72E958A0E9AEE955670D55A31F79D7D09D150CA14EC5204CD9A85ACA00906",
		INIT_1A => x"3C31B9881C3A7D2A057373DBCFF9DBBB1CBF9159BE73FDEAF4FBEF21A37C1EE3",
		INIT_1B => x"0C336ACBD57CC4AAE28AD12B0D33A4E73425E4FB5ACA63FA946DA1020744224C",
		INIT_1C => x"DB8768245A16EB5E85F84704330CB8AB010C119BF704A1BDA2FA7CFAB94DBEFB",
		INIT_1D => x"8D16CD68E0EC779E188BDE89C88CC40CD2B98EE5EA2695A509FBB8CBC2C658DA",
		INIT_1E => x"155D4BCF20A36F40E8268D601634D266C4635A9B203DEB4B27000C588D9EA948",
		INIT_1F => x"CB7CFF4C454E16146B168485524D6C86273571E1648ECADD0DA18E0EC374E238",
		INIT_20 => x"B90D9A0845E025F3B3AECA526A595A7F71BA0D1FE84B28B4054DC05033C2DCC1",
		INIT_21 => x"209A694EDFC866C3F634AB5FB76493950FAFAA82EC27665D1948AB5239736C08",
		INIT_22 => x"5C76B7EA4749F63D594E1DFCBDC8BE14DEC4FB6B4A7F4A5B7BC33A8E13145C27",
		INIT_23 => x"922E8DD7B39B4784C2FFB74D4B98E773C4B69DE1401F700DA13C93AF6764AE06",
		INIT_24 => x"CDBFE0585E940E0771AB0958C4046C052E63E10012A484683DF1CDD7A5D0DF2A",
		INIT_25 => x"F063EE6609945CD61CAC0B8FC17E7A42DDC34A29FE3C86D724F26EE914A3916B",
		INIT_26 => x"0009A5AEAD8B9280934AEC1DDDE49256725EE1C85F6D2EA5E98D27F17621A11F",
		INIT_27 => x"40DCB9FB2E72F9379F6ABCAD98B68DDE8CF726240DCD53D422B9974372415CA2",
		INIT_28 => x"BE8D62EC661F1402122DD62A932141D4B56029DB9A7D2D2437E34CC8572BF7E5",
		INIT_29 => x"11AB90C3F4ED07FD899BD1D82BFA04FADE1532FD8F56F968FEA6949C4F7548DC",
		INIT_2A => x"DE67528D7C3AF34BC3572F7871C952C0916052CAA4471C958C827BA4FEC7AA0B",
		INIT_2B => x"7302713DE8AF0670FDD1078B09749FA553361303E14B73E97A977BAEA996FEFF",
		INIT_2C => x"495853845879EEA0C4DAF10BE8C5E594764FA55196FA8A9F55918A199F196308",
		INIT_2D => x"15057DE4E77054A24AACE86D93D53576619DC943B94228E7C2C0BD9D3D43C56A",
		INIT_2E => x"886914323D3305D77373209B073D14D3DA9385D4F8E7832C02486892E5E6BD03",
		INIT_2F => x"95F02FC83FC4345A631AE3286DD6ED480440A6D338E1C0D5599F97AB510E4B88",
		INIT_30 => x"435383BE91C149262EAF5EC50F34E031497F21DD59138AD0FE18BAFC183D2A62",
		INIT_31 => x"F2E4835C1E95C1078193E94CF89460E53FFDFB9DEF723D25E28ABB36677AD638",
		INIT_32 => x"499DE4C6727C5D49285850DB07F6DB573E5132F6FA72B25829BCAE8E7F81B4B3",
		INIT_33 => x"1FB1864BCC1D91B43E925947F1624443E8AB4A484B4BDD6D19386F9B157F9764",
		INIT_34 => x"3A9037D8BCDA90F07DD450B1D7A5FD1ADB2B5AB71D7CC796F8454215539FA071",
		INIT_35 => x"CB5EB7F45DF6EA70CB8BBC45E558064AC7195FA0FC52C8BECA9934936E0791EE",
		INIT_36 => x"1C1044CF8D54AEC09561344F9668466EE900665A511149E00E45E175301309A3",
		INIT_37 => x"47AD5FAE1A5005CFFD5B30D77CAF5533371DE662C77273594DA44FC726672265",
		INIT_38 => x"CFF9CEF83CE4FCF499BC212962BABCB52EA43CD7DBA6186FF619802A23107D22",
		INIT_39 => x"A6E3AFFCFBDB457C6C1908A0C367E1B5D9A5BF439EA8E236D49805B4A54788E4",
		INIT_3A => x"D888044A58E6E650AD6B91780DF299B0A3BD703866D3A5A02A4CE2B85497D2AE",
		INIT_3B => x"102B734536311A4AC9125B887F081F3900A17F989A4FC9D923AFDE0FCA130B2E",
		INIT_3C => x"50EBC11C0A7F0428057DD9E59375867DEC99D1DCC1BE6A35CEE0B1D5AEA376E6",
		INIT_3D => x"761AEE5105557857FC8A534F875AD0B03FB7E3E49DF8A98DD2DC48D5114EE0D9",
		INIT_3E => x"6756891676285CEF619C775626C1B205E77EC9943C28711BD93B768AAE6702F4",
		INIT_3F => x"F15917D9EF183AC1EE5A613D5F23831C65DBF2F001577D1424F5691294AB7CAD"
	)port map (
		DO   => doutout,			-- Port 16-bit Data Output
		DOP  => open,				-- Port 2-bit Parity Output
		ADDR => addrin,				-- Port 10-bit Address Input
		CLK  => clkin, 				-- Port Clock
		DI   => (others => '0'),	-- Port 16-bit Data Input
		DIP  => (others => '0'),	-- Port 2-bit parity Input
		EN   => '1',				-- Port RAM Enable Input
		SSR  => '0',				-- Port Synchronous Set/Reset Input
		WE   => '0'					-- Port Write Enable Input
	);
	-- End of FRAME0003_RAMB03 instantiation

end FRAME0003_A3;