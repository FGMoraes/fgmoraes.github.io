--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
--	Grupo de Apoio ao Projeto de Hardware  - GAPH
--	Projeto X10GiGA - FINEP/PUCRS/TERACOM
--
--	M�dulo:	Mem�ria - Gerador de Frames - Prototipa��o
--	Autor:	Jeferson Camargo de Oliveira
--
-- 	FRAME:	0000
-- 	RAMB:	02
-- 	CONJ:	B
--
--	M�dulo gerado em 17 de July de 2008 �s 16h55min pelo
--	programa gerador de frames OTN do projeto X10GiGA.
--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

----Pragma translate_off
library unisim ;
use unisim.vcomponents.all ;
----Pragma translate_on

entity FRAME0000_B2 is
port(
		addr	: in  std_logic_vector(9 downto 0);	-- Barramento de endere�os da porta
		clk		: in  std_logic;					-- Entrada de clock para a porta
		dout	: out std_logic_vector(15 downto 0)	-- Sa�da de dados da porta
	);
end FRAME0000_B2;

architecture FRAME0000_B2 of FRAME0000_B2 is

	signal addrin	: std_logic_vector(9 downto 0);
	signal clkin	: std_logic;
	signal doutout	: std_logic_vector(15 downto 0);

	component RAMB16_S18 is
	generic(
		WRITE_MODE : string;
		INIT_00,INIT_01,INIT_02,INIT_03,INIT_04,INIT_05,INIT_06,INIT_07,
		INIT_08,INIT_09,INIT_0A,INIT_0B,INIT_0C,INIT_0D,INIT_0E,INIT_0F,
		INIT_10,INIT_11,INIT_12,INIT_13,INIT_14,INIT_15,INIT_16,INIT_17,
		INIT_18,INIT_19,INIT_1A,INIT_1B,INIT_1C,INIT_1D,INIT_1E,INIT_1F,
		INIT_20,INIT_21,INIT_22,INIT_23,INIT_24,INIT_25,INIT_26,INIT_27,
		INIT_28,INIT_29,INIT_2A,INIT_2B,INIT_2C,INIT_2D,INIT_2E,INIT_2F,
		INIT_30,INIT_31,INIT_32,INIT_33,INIT_34,INIT_35,INIT_36,INIT_37,
		INIT_38,INIT_39,INIT_3A,INIT_3B,INIT_3C,INIT_3D,INIT_3E,INIT_3F : bit_vector
	);
	port(
		DO   : out std_logic_vector(15 downto 0);	-- Port 16-bit Data Output
		DOP  : out std_logic_vector(1  downto 0);	-- Port 2-bit Parity Output
		ADDR : in  std_logic_vector(9  downto 0); 	-- Port 10-bit Address Input
		CLK  : in  std_logic;			 			-- Port Clock
		DI   : in  std_logic_vector(15 downto 0); 	-- Port 16-bit Data Input
		DIP  : in  std_logic_vector(1  downto 0); 	-- Port 2-bit parity Input
		EN   : in  std_logic;			 			-- Port RAM Enable Input
		SSR  : in  std_logic;			 			-- Port Synchronous Set/Reset Input
		WE   : in  std_logic			 			-- Port Write Enable Input
	);
	end component;

begin

	addrin <= addr;
	clkin  <= clk;
	dout   <= doutout;

	-- FRAME0000_RAMB06 instantiation
	FRAME0000_RAMB06 : RAMB16_S18
	generic map (

		-- The following generics are only necessary if you wish to change the default behavior.
		WRITE_MODE => "NO_CHANGE", 	-- WRITE_FIRST, READ_FIRST or NO_CHANGE

		-- The following generic INIT_xx declarations are only necessary
		-- if you wish to change the initial contents of the RAM to anything
		-- other than all zero's.
		INIT_00 => x"4BEE9847560F7C825BDB7ECEA6846859D85C5532B20B90C12D90D3BB6811E741",
		INIT_01 => x"EA35DD7CC9195CC84E06F4858BE0FAA7EB41250C0B79A7A5B07BE58079707DCE",
		INIT_02 => x"9A9DB96BACC616E06D67E21B159D422C3DD3FAD01B6B1BB57A8744751610A70E",
		INIT_03 => x"C6E4E7EC77B47B472997214A60B826788054E10B811A35328C338DDAF900E83F",
		INIT_04 => x"D848D06515CD2B5B48585E2651100D87E2B36D7A4EA4E27CB4F44E5037096B8C",
		INIT_05 => x"3F753E4237B22E82AB5D896F6CD4EFA1BAD0F0DC95141F1FC2513B41F0E7A78A",
		INIT_06 => x"79E82CBC64A1CB8CC067A311F3DBA7F51B87E01CED7127C51D7CD893D5F35235",
		INIT_07 => x"4E305245CD75CFEAA0BA9B4F871F6DC3C072F5446BE10302A2B41FA92BC9413A",
		INIT_08 => x"151280AE972DCE2251F47CC1A1C8FE80B1F89864CB6DA6F2D0EE712DEBB56E02",
		INIT_09 => x"013F3CAEC8AA0C1212A63F546525019E880C738403026E7BE2FDA241A44662A4",
		INIT_0A => x"44795F8485FDDC4902C8EF111E05D4B19E81D89770ECE6B14C0769794A91B2D6",
		INIT_0B => x"CEE5726AE1B8A8B0FC23CF9E2A472B030A3C0B91D089FBBAC42EE25699A6C13D",
		INIT_0C => x"F1B433740A76F4B1CA6D1A9BA047D9B8EEECE36C45FA7CF28F2AE4FEBB1DC950",
		INIT_0D => x"5CC9345148B63EFD10177BC78E4C345A05D51290752A84A3DD817B5C2F2257E1",
		INIT_0E => x"B6F274116209247977EA3822B760EEBB2C0EDCEF3B36156EBDF4290363419C8D",
		INIT_0F => x"EFACAD7C2C08E51CC2B96347C930833C3EF8EC1BF14FF8B1A59A7B82F2DCFB32",
		INIT_10 => x"A0EE7646E4E77DAF8CCE808F86873ECA3CF61527D3ADE8D9CC15EC663945FC49",
		INIT_11 => x"060DDDAE7112C4341190DD6636D09C543E80A2325EF4AF4536FF434DC4FFB154",
		INIT_12 => x"D707E122B182CFD723B5C259DB927A176AAFE8635C1AC100467AF7181406801C",
		INIT_13 => x"AD180F4ADB4B67DAB5D560FB856EADEC344187D67ADF5C3EA1162F9F4DF8A423",
		INIT_14 => x"E5505354B7E7419C4D9A2536DCA655724D1AFA9C8979C446B0E81EEC94CB846A",
		INIT_15 => x"264BF8FB8FFF4BA9F0BC0B36667E49D4774FE66B56B48DB8F39C14D7EF49BD92",
		INIT_16 => x"4BE77F96A0D455BDE5667D16D7E5EAEBA4FC57AA79903B26135EAD30AF96F766",
		INIT_17 => x"201EF13DC47C3985D220C2E1E71A2D17845B788D838F184337CD6D7512BCD3F4",
		INIT_18 => x"029AF5B6DDE9B8BDCE181178E59CAEEB9296EBCCB2A37171BCE2CE7FBA8E9C50",
		INIT_19 => x"8A922630F9959EC238086D7AD300D19552ED2AE450F5512B8050CD3BCAF3708D",
		INIT_1A => x"844FAFAA45FE0E046E7ACC2FD7402E211856E4D782A320E2A35D0FEC6D4E5AF4",
		INIT_1B => x"8FAF04EF3ED58C388E083E8AE8E93A5ADB115585B953D991492FABDA24951D74",
		INIT_1C => x"7B6419862F7F44FA69E06B6B9A460CB739B2C42FD3C70D3DF8E83D5EB2273077",
		INIT_1D => x"4A367DE7DDD6D2A1E19C75793462825EB7BA00C5630500224390C2F677233425",
		INIT_1E => x"F6963D05182945878004FFD9526697A996A071EF3D85155121727F35322BA96C",
		INIT_1F => x"210C191183150EC472BFB4EE3997DACFCDEB7E92A0FFA00B4A9413D74AC71702",
		INIT_20 => x"78D1502C527FC04C516703B88934351592A2327A2F39BD714797F78493E22052",
		INIT_21 => x"C9961C8622AE70C85AAE486BDC1D38A612172A629B3E8DBB6366A04FA8D62646",
		INIT_22 => x"6236471665C1018A9C046A89925702FE9F84986A49ECC9D020A2E36B8DA5CAE0",
		INIT_23 => x"0C3008246D4351297AB6C8D805C456259454B6F70F2C437B3A94171E7B487053",
		INIT_24 => x"83FC5BD88C0C8BA733DE41AD5E06117A94884C7156AA423D313535ABC4DD7B2B",
		INIT_25 => x"D44B735983F36B49B0A04232DE7F3CEDDE0D2B24CD51B02B970FFD3A36800142",
		INIT_26 => x"3331CC4394A5A68EE4070A566241C109543C472AE9E7FF866B11580410DB7A01",
		INIT_27 => x"F63DF6DA53C2DD564464F2CBC2DFF1F33091E771628642824644011823351C1A",
		INIT_28 => x"31E8CFE34846FA4EE5B16C7DD6516CB5F71EEC45CC5A7428F863E904D1F997C9",
		INIT_29 => x"A60C4A0B0EF9D6D9542CF412FE611A18D140276BA64FFF1F39A607A4C904754E",
		INIT_2A => x"7953DC788EF71813A628DBF6D1F2230A0FB640B28A025A6D38319E76B39B755B",
		INIT_2B => x"F4853C1C44D15CA82A2EC626B80A22806A8C5BB32B6BD3A74BC851361DC63BB1",
		INIT_2C => x"24BB75F61622D6E57E880D0A9B1F29E428ECD06BBE6B0F7D50A0F0C78711E204",
		INIT_2D => x"6C14A52215A0A0F5BF829C6F8B442319CE6E535149BDFE366DAC2B03A912172A",
		INIT_2E => x"74B9AC479775AFB54FA4021DDBD51C4881EF56FE8D7663B86251106A61D063D8",
		INIT_2F => x"E7AB173D33BD6F79F8A5469A998A8E3C74B04F3CA406C88177EE72035CEC60F8",
		INIT_30 => x"E811BCB84DEE57CBF8C16F99F314638E379FE53645FA3CBC22B067D08BA655CC",
		INIT_31 => x"02432FD7DA5C4002E738FD97A04379F5EEE3459A8F572EE026F076B75601BE35",
		INIT_32 => x"9680B94E09B0F9801756295CAEBDB970C4F7B6F6A486FD8ADC92CA72E6990427",
		INIT_33 => x"26BD1F2E9CF68DE66461620A6B4E37375AA3047D5CC8323E4648469CF8FA4659",
		INIT_34 => x"92207D8388A0F2F1AB3495FFBBC944DD0A756FBAB9891806CDFFDE9EFE1C00DB",
		INIT_35 => x"339324B19FB72AD0FA37072814754D289DFFB28ABDFFF81E8356F9C4E57307A1",
		INIT_36 => x"258D325AF944203F356980BC202D55A10583967FD1D1FADB06C25377C065DFF5",
		INIT_37 => x"612B6B74A10DABBF1664D40D040A5C86E98246F7CF9F1DF30A69E7C77E32FCB2",
		INIT_38 => x"605677648A128F2FBE8C652E6E29084D2AE51432636375F4F521308CC8616A11",
		INIT_39 => x"CD5839720B1CAA2CC62B318E48261899D6BDDCB77BD8B62B793FBF8A38EB62C0",
		INIT_3A => x"9393F7B92C5F5A04135B302A7EDDDC4A739818C6D01D2639A3DC22234E633D63",
		INIT_3B => x"0E9FE064AEE78C801661912E8A164CEA1C4C45E0078E3BD3893C7D213D7BD701",
		INIT_3C => x"35B26CDAE4C374D7D400D81C4742F52EFA15AFC2AD2EAFEE80A0D950A852AC2A",
		INIT_3D => x"29AE90446529845C8179317ABCC8CAC452CCBAF22BAA2005A2EB6C03680FC774",
		INIT_3E => x"2443F654DDD65657D935396DA0572947B93AB5C9C8D8B427B0515D5781083D41",
		INIT_3F => x"111111111111111111111111111111113F3DF54CD33DD14660D1A99E45C9B8B5"
	)port map (
		DO   => doutout,			-- Port 16-bit Data Output
		DOP  => open,				-- Port 2-bit Parity Output
		ADDR => addrin,				-- Port 10-bit Address Input
		CLK  => clkin, 				-- Port Clock
		DI   => (others => '0'),	-- Port 16-bit Data Input
		DIP  => (others => '0'),	-- Port 2-bit parity Input
		EN   => '1',				-- Port RAM Enable Input
		SSR  => '0',				-- Port Synchronous Set/Reset Input
		WE   => '0'					-- Port Write Enable Input
	);
	-- End of FRAME0000_RAMB06 instantiation

end FRAME0000_B2;