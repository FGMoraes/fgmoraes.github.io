--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
--	Grupo de Apoio ao Projeto de Hardware  - GAPH
--	Projeto X10GiGA - FINEP/PUCRS/TERACOM
--
--	M�dulo:	Mem�ria - Gerador de Frames - Prototipa��o
--	Autor:	Jeferson Camargo de Oliveira
--
-- 	FRAME:	0002
-- 	RAMB:	00
-- 	CONJ:	B
--
--	M�dulo gerado em 17 de July de 2008 �s 16h55min pelo
--	programa gerador de frames OTN do projeto X10GiGA.
--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

----Pragma translate_off
library unisim ;
use unisim.vcomponents.all ;
----Pragma translate_on

entity FRAME0002_B0 is
port(
		addr	: in  std_logic_vector(9 downto 0);	-- Barramento de endere�os da porta
		clk		: in  std_logic;					-- Entrada de clock para a porta
		dout	: out std_logic_vector(15 downto 0)	-- Sa�da de dados da porta
	);
end FRAME0002_B0;

architecture FRAME0002_B0 of FRAME0002_B0 is

	signal addrin	: std_logic_vector(9 downto 0);
	signal clkin	: std_logic;
	signal doutout	: std_logic_vector(15 downto 0);

	component RAMB16_S18 is
	generic(
		WRITE_MODE : string;
		INIT_00,INIT_01,INIT_02,INIT_03,INIT_04,INIT_05,INIT_06,INIT_07,
		INIT_08,INIT_09,INIT_0A,INIT_0B,INIT_0C,INIT_0D,INIT_0E,INIT_0F,
		INIT_10,INIT_11,INIT_12,INIT_13,INIT_14,INIT_15,INIT_16,INIT_17,
		INIT_18,INIT_19,INIT_1A,INIT_1B,INIT_1C,INIT_1D,INIT_1E,INIT_1F,
		INIT_20,INIT_21,INIT_22,INIT_23,INIT_24,INIT_25,INIT_26,INIT_27,
		INIT_28,INIT_29,INIT_2A,INIT_2B,INIT_2C,INIT_2D,INIT_2E,INIT_2F,
		INIT_30,INIT_31,INIT_32,INIT_33,INIT_34,INIT_35,INIT_36,INIT_37,
		INIT_38,INIT_39,INIT_3A,INIT_3B,INIT_3C,INIT_3D,INIT_3E,INIT_3F : bit_vector
	);
	port(
		DO   : out std_logic_vector(15 downto 0);	-- Port 16-bit Data Output
		DOP  : out std_logic_vector(1  downto 0);	-- Port 2-bit Parity Output
		ADDR : in  std_logic_vector(9  downto 0); 	-- Port 10-bit Address Input
		CLK  : in  std_logic;			 			-- Port Clock
		DI   : in  std_logic_vector(15 downto 0); 	-- Port 16-bit Data Input
		DIP  : in  std_logic_vector(1  downto 0); 	-- Port 2-bit parity Input
		EN   : in  std_logic;			 			-- Port RAM Enable Input
		SSR  : in  std_logic;			 			-- Port Synchronous Set/Reset Input
		WE   : in  std_logic			 			-- Port Write Enable Input
	);
	end component;

begin

	addrin <= addr;
	clkin  <= clk;
	dout   <= doutout;

	-- FRAME0002_RAMB04 instantiation
	FRAME0002_RAMB04 : RAMB16_S18
	generic map (

		-- The following generics are only necessary if you wish to change the default behavior.
		WRITE_MODE => "NO_CHANGE", 	-- WRITE_FIRST, READ_FIRST or NO_CHANGE

		-- The following generic INIT_xx declarations are only necessary
		-- if you wish to change the initial contents of the RAM to anything
		-- other than all zero's.
		INIT_00 => x"D3D8BFBBBBA26B888FF179CE2B82D288DFDE995933D00A4752D1B856C1AD6C9B",
		INIT_01 => x"B6670937C84BFFBC2A36F7A3127477E92BD8E1EC4C853F337B048FA0859C23B4",
		INIT_02 => x"D24DFF92B2AD37E66550BCDC64BF0B15A700B81D0E0338EDC4B942E57CE59FE1",
		INIT_03 => x"13940F6ABD462622F0075FAE1E810D7F09BB330BBC79D6641AA71D1765CEA805",
		INIT_04 => x"41107709053A4DA3CCA7342058A373116D6D2BFF3B23523CF729C345B7335566",
		INIT_05 => x"76D7AE863E56DE8FCC8A2347244582B424C5E6ECFBD4470A90180B7134C0517D",
		INIT_06 => x"919260EACC662188A777F44E9956D748B85E249DF0370AC0311754B1B9F3A24B",
		INIT_07 => x"245B16F020671902D164E4BFBDEDA82865DE15EF2ABBC34BBC5F34B4FCC685CF",
		INIT_08 => x"C52610DB46A66D9678704028FD2D956536654B48575CCEC2A35EE38DDF8DD757",
		INIT_09 => x"489124A863EF27466E8A314D0474B46CF527486FF1B25BEF6602E7F8C004D999",
		INIT_0A => x"7D452DE6F189737580F69081B263E3D48F98BE511A30015C1927D34ED6387FCB",
		INIT_0B => x"67D2E8C02CECE8392959BD62704D8DB33E69779C38331EFDB3B32E7362267781",
		INIT_0C => x"07415E93455C0F66AAAAFD5E81D42D976E94C4B04C3FB22B028C951EA994FDBD",
		INIT_0D => x"134D7AF333BD7B1D235087AB707A6BB714036F9A3D73E012C2DF070A69F16190",
		INIT_0E => x"7DEBD551FB12372E651114D12CFE57522ED724147F8E692592FC3EFD9DAA96AC",
		INIT_0F => x"0A5C934C41977975576FE7557F7EB7393839521AA5ABF335173C67D45E1880CE",
		INIT_10 => x"D20E5CFD8F3075C4C84965ECDD259C1F921F4FDDA75AEE0B889E785D9593D10C",
		INIT_11 => x"97C24C9DBB05E086F24772F56F4CAB6075A0A5BFBCC4C018D6C54EC62D512BF7",
		INIT_12 => x"CC2C5EE2CCBB4250D17C423FE37A1C0C940A7F89DB356125B4185F9DCCD39E89",
		INIT_13 => x"EF45EDB27B015C8F968280F7820E74A05F2702AE38F1722968E2DC476150ABB7",
		INIT_14 => x"4080E8DDB6002E5B924B073F18B1A92C192A2469CF897C281B75A96566071420",
		INIT_15 => x"EB5CD249C6BA867FB506E5CB6EC8FC0BA529C1B59AD8728DABDF316B2D6D957D",
		INIT_16 => x"39EFB784AC27FF907F32AED0CDFD0C7FCF6521C523723C6659E8CE559B21A822",
		INIT_17 => x"7C451E04536B8D166060FAC7D214AA762D950DEDDC2B5F436924C3CFE867C821",
		INIT_18 => x"C4AB31D074A9F94CA242CDA13EAB65D7A30EA7AFA9008D217A8D7B1E02D227D7",
		INIT_19 => x"0C6A9E190A3611FB1D67FB4308D6FFDE83559560F8A4071846FE25868A9E2C9D",
		INIT_1A => x"1081A8CF22D4784EA45B1D98FE026E20D660C923C2446673654B7ED2A6C16D5A",
		INIT_1B => x"8987A9040AF60A03CE194D10A2A10B30C5BE384DBF1E6944B6444637B2FACA66",
		INIT_1C => x"597075B3BE7EC164C77A1E3D81BAE023CE46A659D96F921EB74C290BABDF99CA",
		INIT_1D => x"738F7C0575A830CE47474EDC41143BA3D651EABF3CEF384C7D4E48BC4A5B80AA",
		INIT_1E => x"215CB98A51A4362B164443716C5A13483D7BF885638360103F8DD9384B0AC111",
		INIT_1F => x"9AD2103B2BE2012BDB7446E1BE404FCCB4DAAB7F5D6DA0554082F42CCA073B0A",
		INIT_20 => x"25733C69C649B4E3EAB80DF0C1EF23B6233CD1093A9713C752D164EB28CA4C20",
		INIT_21 => x"A622020405290ECFF20A2E0976813DF3141E9A71733F046DC517A9A29AD4595C",
		INIT_22 => x"5686745F045DC8986E3A6252012B97051D6280EFB51CD4C516F271FC4BAC483D",
		INIT_23 => x"80BB9048389B24AC19CB571C7604B19CD6A035CC08238629A99E33CF4759C11B",
		INIT_24 => x"64F133667BD202BE02961E439B557B68E9B078FD7B62D460970770F920C71B48",
		INIT_25 => x"602BF24CBCCAB154079841878D4BFFA64AFB917655DD86EFB5382108BE99453C",
		INIT_26 => x"FF0A794B2593B489C1B986E5C753059AD51B15102F5CDC3D0DA339166CEFFEBA",
		INIT_27 => x"B86A94448A25426454415065AE50C55AFEAC0A8414E310062CD56754DAD2E2B4",
		INIT_28 => x"14C691AF9E962BFBE34507863127F23181D332EFCC47782A27DD98CA61566484",
		INIT_29 => x"0928A6D60F79111B188A7024CD2491D99EEAF95629803D303898B97FC9E45477",
		INIT_2A => x"6583D7AB1144D11639E997D757D0D0ECC3C3379C0C90E7D18BDFF32E918A94F1",
		INIT_2B => x"DF56AA4B5E5541C8AB068818954F660C2E412564015D17FC5431D7822A3E8DA4",
		INIT_2C => x"2524CA9E66687A0B33F0729E0FC630A92B16F45B23AC12C2ABDC67F87A43ED9D",
		INIT_2D => x"F9A6C3706E24779C8FDF83C3A0EBDDC0EB37194FEEEE838C23A3F1092C1F6857",
		INIT_2E => x"69DE4FA34FCC3F2F1D2DE136D8A2FBC894361B1E852971D91BFC8C4FB7335510",
		INIT_2F => x"56F8F83ACFBB8F6372B830F0307D3C797C9AC2F47497D4CDB3DA74204180A9F8",
		INIT_30 => x"88DA14F335319C1DF55392A6052F8D00E84A1E0D5029486EC06BD2726215E648",
		INIT_31 => x"1A50574C7EBBEFAB2B3D8C5DBB7D99208608C210754E559860105CC38E4CDE29",
		INIT_32 => x"9FDA4808D769C92598A8F0A8C9661095870877025A100EF7543DF439F391F48E",
		INIT_33 => x"69C61C9385ECB278F3CCF1EE3ABFADCB0873FC032A16CA097B7FE4F943577AA8",
		INIT_34 => x"1937AD90B41C22351EB8A542171E21CE67527F61EF028E545F0D52898B981E1F",
		INIT_35 => x"E54B47977B7E9CD0688C73CFB35725B67C38D30B1BAFBFE2DC023C588DD90845",
		INIT_36 => x"5DC3105FEA305DDD4337E5AA6ED92040426E1E33CCCB1D3288CB708071CC23F1",
		INIT_37 => x"95750F6294C0A0C21B74A7B09AAE8F6ED114AB64830EFD53B4BF510A4B4D1CA1",
		INIT_38 => x"066498A932704A6C1BBEF636AE8567AE8283AB8020DD2A28BF86548E3CEA1BFA",
		INIT_39 => x"311CC794C850F8A46834440B12794609F7101BBF25D98C10F31AFBA330BAA56C",
		INIT_3A => x"72FBF3D9066AFF6D772687B0CD82DFD988830AB9B15E2A92AB237A371F741710",
		INIT_3B => x"6644BE7E675078C0AEBF2DB661185C892A2145776EC13DCB18C6BCA374BBEE15",
		INIT_3C => x"B32480F650DFB8A7A14F6EA5B66E93888A76B36DAB79732304EB3C900FCB4B0F",
		INIT_3D => x"25ADD2C9426668CF1D67CC3FB38DA1512C9F79D95885921865E9DB2D2D6AA7C5",
		INIT_3E => x"1977D9D18B2E2F8517177A4C985DAB75EE3AEEBA4E0CCE17FB3658B8B2D4D6D5",
		INIT_3F => x"11111111111111111111111111111111422E7F845A7DE91809DAD0EFBF893CDF"
	)port map (
		DO   => doutout,			-- Port 16-bit Data Output
		DOP  => open,				-- Port 2-bit Parity Output
		ADDR => addrin,				-- Port 10-bit Address Input
		CLK  => clkin, 				-- Port Clock
		DI   => (others => '0'),	-- Port 16-bit Data Input
		DIP  => (others => '0'),	-- Port 2-bit parity Input
		EN   => '1',				-- Port RAM Enable Input
		SSR  => '0',				-- Port Synchronous Set/Reset Input
		WE   => '0'					-- Port Write Enable Input
	);
	-- End of FRAME0002_RAMB04 instantiation

end FRAME0002_B0;