--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
--	Grupo de Apoio ao Projeto de Hardware  - GAPH
--	Projeto X10GiGA - FINEP/PUCRS/TERACOM
--
--	M�dulo:	Mem�ria - Gerador de Frames - Prototipa��o
--	Autor:	Jeferson Camargo de Oliveira
--
-- 	FRAME:	0000
-- 	RAMB:	03
-- 	CONJ:	B
--
--	M�dulo gerado em 17 de July de 2008 �s 16h55min pelo
--	programa gerador de frames OTN do projeto X10GiGA.
--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

----Pragma translate_off
library unisim ;
use unisim.vcomponents.all ;
----Pragma translate_on

entity FRAME0000_B3 is
port(
		addr	: in  std_logic_vector(9 downto 0);	-- Barramento de endere�os da porta
		clk		: in  std_logic;					-- Entrada de clock para a porta
		dout	: out std_logic_vector(15 downto 0)	-- Sa�da de dados da porta
	);
end FRAME0000_B3;

architecture FRAME0000_B3 of FRAME0000_B3 is

	signal addrin	: std_logic_vector(9 downto 0);
	signal clkin	: std_logic;
	signal doutout	: std_logic_vector(15 downto 0);

	component RAMB16_S18 is
	generic(
		WRITE_MODE : string;
		INIT_00,INIT_01,INIT_02,INIT_03,INIT_04,INIT_05,INIT_06,INIT_07,
		INIT_08,INIT_09,INIT_0A,INIT_0B,INIT_0C,INIT_0D,INIT_0E,INIT_0F,
		INIT_10,INIT_11,INIT_12,INIT_13,INIT_14,INIT_15,INIT_16,INIT_17,
		INIT_18,INIT_19,INIT_1A,INIT_1B,INIT_1C,INIT_1D,INIT_1E,INIT_1F,
		INIT_20,INIT_21,INIT_22,INIT_23,INIT_24,INIT_25,INIT_26,INIT_27,
		INIT_28,INIT_29,INIT_2A,INIT_2B,INIT_2C,INIT_2D,INIT_2E,INIT_2F,
		INIT_30,INIT_31,INIT_32,INIT_33,INIT_34,INIT_35,INIT_36,INIT_37,
		INIT_38,INIT_39,INIT_3A,INIT_3B,INIT_3C,INIT_3D,INIT_3E,INIT_3F : bit_vector
	);
	port(
		DO   : out std_logic_vector(15 downto 0);	-- Port 16-bit Data Output
		DOP  : out std_logic_vector(1  downto 0);	-- Port 2-bit Parity Output
		ADDR : in  std_logic_vector(9  downto 0); 	-- Port 10-bit Address Input
		CLK  : in  std_logic;			 			-- Port Clock
		DI   : in  std_logic_vector(15 downto 0); 	-- Port 16-bit Data Input
		DIP  : in  std_logic_vector(1  downto 0); 	-- Port 2-bit parity Input
		EN   : in  std_logic;			 			-- Port RAM Enable Input
		SSR  : in  std_logic;			 			-- Port Synchronous Set/Reset Input
		WE   : in  std_logic			 			-- Port Write Enable Input
	);
	end component;

begin

	addrin <= addr;
	clkin  <= clk;
	dout   <= doutout;

	-- FRAME0000_RAMB07 instantiation
	FRAME0000_RAMB07 : RAMB16_S18
	generic map (

		-- The following generics are only necessary if you wish to change the default behavior.
		WRITE_MODE => "NO_CHANGE", 	-- WRITE_FIRST, READ_FIRST or NO_CHANGE

		-- The following generic INIT_xx declarations are only necessary
		-- if you wish to change the initial contents of the RAM to anything
		-- other than all zero's.
		INIT_00 => x"A88EB8FD636D0AD78E67128938BBC9F71F4535E7FDBFF83936F91A247498B0D2",
		INIT_01 => x"CCF80F647311625FDC4C3F8532711E2B844D611332DEE721D22EFA0D06D0E977",
		INIT_02 => x"6816A1C1DFF0EBD3EEB98C2CD7C2FAB10C785CA2C37AD247C684E5E9E24C88EF",
		INIT_03 => x"39688D2C0D71CA6962DA5D2ACFBA4E2B633EFCA862CA1030DDBFFCD6029411A4",
		INIT_04 => x"65A16E7268A52AD83E0BDC063586A77012ED744B866A79D21154070597584D00",
		INIT_05 => x"E8D4C6FC2D505845F333B20FC0F1BE0F6E6D2CC2232A676CC51B87AFCB21EA6E",
		INIT_06 => x"283BCB1C3F4BA4BEAB75BFAAFF42B2929FA60AB7F52FC868725BCD73E8C666A8",
		INIT_07 => x"4F6CFBA64C35294872518D71DC9A789806073548F4FA6E1BF698CEB7DECD5329",
		INIT_08 => x"1E19FD0139BDFE0BF9364B4A9EDE5A7DCDC7A8D1E68348D378CE0D71032F4DDE",
		INIT_09 => x"30999EE04B1453229B39C17CE6850A387FB040644A9DE6EC3D57882A324D4A74",
		INIT_0A => x"5809E95164F19F03C7A8C8D7BA5E19EFCCC6E466DFC73D0B454FBF27618D237B",
		INIT_0B => x"9C78824093FFA9898AF4256230164D72595CED01A32BE0F31AE5E10A39909811",
		INIT_0C => x"E0DD2CDEEA985D996023788568EA3A3D2A4B14F7A9AF34EBD26B6C01F55A65FF",
		INIT_0D => x"024993201998318EDBF40E444B2833E6C1BE1E3BFA744352F7CA993EC6ED596D",
		INIT_0E => x"0BB9DB395AA61DE0B2AE4BED88F9918B2F05D78AD58D0C5A3A64B6D5EEDDB61D",
		INIT_0F => x"3825BF3600D4DC99AEC0D69635F8365AE0BC4364E2A8F0D516692AB0040AC500",
		INIT_10 => x"E38243AB0C9B0ECC98096734D522361E142C0A41F94C25DDB02177ECFFB83C43",
		INIT_11 => x"A930A1549A5BEFB824453FA9EA7B7499ED7D4E71B59D1F20CF1C851B82BE615F",
		INIT_12 => x"B26DB9AFD358948FD2704B9BDAFD715DE715B2A0A94D9D287F730E537ED468D5",
		INIT_13 => x"FAAB332A3F2FF0D677BA21554B988BE97A8724FEB60228A996F3557190F199BE",
		INIT_14 => x"AEC04B3D7505BDB9B8DC152406AF13681F80F7132C9D84BCFB1397A5D6A69F14",
		INIT_15 => x"A685D42046BD54DE02E5B848CB97B63E8B930D6B7D8D8BAB14A527E19A988D6F",
		INIT_16 => x"561F09BE8F78044D2CB58F565813541907C249391AB75DF7E4D3C9001C630D2C",
		INIT_17 => x"FCAB967A36FA729A90DD9DAD85ED64F03A2DF28F7EC15CD96FAC575A9ECBB092",
		INIT_18 => x"600D32D1FA328881E3DE9DF49F0AB3133BE8DE1612D02632D4DC752D941A827B",
		INIT_19 => x"EA10E6315333964C0C927FB1B17A61645F52F0D639DF563B4E0B5E89E4B5BE0C",
		INIT_1A => x"E54D25D343BE0FF31CF7A10A5524D9B5D8F4E9FCA5CE2120EBAFC041EF30E821",
		INIT_1B => x"7B31B9ED95669667B1695964760978B13FD0276FE7F48485D1FC4BF809091255",
		INIT_1C => x"537B222ABD16BC0D8E05840A0E324F8171ACBDC28E43339104D5016FE97F27F1",
		INIT_1D => x"B0380988C9EA36502C0A5990A8392AC94CE74EA98AA49F22D66107F3A19A29E7",
		INIT_1E => x"AF6F605294C70B1D89DB507035105DAF5F23BFEC902E46F31106ABF8B5B1D6D8",
		INIT_1F => x"4C74EBEEE6E7AE35287C2A7D6CC751BA6ACDEF47141BE076FA6DBF1280EAEB0F",
		INIT_20 => x"FF981E0C71C1604C0B0D8FCDE457D7ADFA5F7E02E361C0F50E387040A64DA81D",
		INIT_21 => x"D2F2B732C6012D2634D073A40F9626B69BCDEBEAC9DCE8CD0AB78DD51D10829B",
		INIT_22 => x"E7BCD7A43600685A19E9491AE6C3AB65E78A98034B78A574D7D5F4741E7EAD8C",
		INIT_23 => x"218BDFFC6943994F6F8574F50796DB55E7E320CCBB7A1DE62EC9DC2739E3FE1E",
		INIT_24 => x"6FDB3F5B928A24DE202D4B65A5FF38F17E6D4D09EE4789693203DD1D8F50E7FF",
		INIT_25 => x"A7F4EB6866542C5D24F74A59BD5C401DA675D81F897D84F53EE0C4C0A6FF036C",
		INIT_26 => x"08F4F33ABD2CB95E92CE5A6DBD9A78F6BA949288834ABE06C96EC6C30FC80000",
		INIT_27 => x"0585E4B2B9916B643D04415C6732780EF2E2AF918B0C61B855F9382EA778C166",
		INIT_28 => x"D30BB86A77C53392F27E9B47E02CDC484DEA1A2C06178975E52E1B262CBAF939",
		INIT_29 => x"678F7BA8143FD7D3658D6D2D357C588F258CD7BBE22D829ED477F1FB5B4D15FB",
		INIT_2A => x"868826913FC34AD2495FE6F64FFDA0F7C84B8E1FB0EAAA80BC91D78416676C49",
		INIT_2B => x"DC855A95E99E92374DFD2760DF8B6DB364BB7E7E2D5079CB6F1CFF81C9FC93D2",
		INIT_2C => x"2F3E6B80B98B91FEF8435CD137383CB7EBA9386B4235DF5D9F0B5D212550AB6C",
		INIT_2D => x"8E43CAD8F6E042EAB71095BAC49BA6306A6F6C42982BF6F89880C20DD3D0F351",
		INIT_2E => x"AD0BF963EBFA76573307DC278FE9B52F43F04ECF79224A2367AB6ED212171812",
		INIT_2F => x"65E15AC5FFD26FAD1E4A4A5B2E8179240D85B51DBC4778EA8D82C000F8DB831B",
		INIT_30 => x"04A514F3FD17A1E81FAFF7D1F7E99386441A02AAE5BA4CB834594E316E7F5836",
		INIT_31 => x"676D31D95D7161C4DBB0EA7497095AB9EC0E182D6177C7434220CA26FA0C1FEF",
		INIT_32 => x"F849EAD2E6214CE52CF501B22B86288AD6AB58EDB3C6CBECD71EBAA69FE5158B",
		INIT_33 => x"8592FB69413A4BDCA92C755F7A6E0FF353B91181E48C973E993C4F80B99082D4",
		INIT_34 => x"BCE29D52E3733916A84CE5782C005B688212BF080E6136EA62AAAA7C70639B8B",
		INIT_35 => x"5929FB99DE3535AD32EC449116E72D1B38AB02491FA3C861E122F66753216573",
		INIT_36 => x"118F4BA3649081602D2C931E46FB9A5170E89F9002AC8070226279FDAAB05F9D",
		INIT_37 => x"A801A912F395FB1ED2C6BA61EC9810B5F89B03F3CA73A88E2759D8614DA37CD1",
		INIT_38 => x"D94B8B36D17591577253E94EFCD829A945C005294E1B683631CDDC34F5418FC1",
		INIT_39 => x"960F47630C34490024791910808B8EF6D359211E861AF7EAD715EE5769A0EEEF",
		INIT_3A => x"F5A556BE750722B667DF5AEC76F3FBA1CF8D46DA7C2B526C47186E2BA667F671",
		INIT_3B => x"15270C393C89707C640D8AC002A4DFBECFAA2D833EA823563D6F6E9DDB3F2344",
		INIT_3C => x"79F3AD1304ABCD7CD454DF90E88C38C987D39007713F2DFC2A88215EAD1BA194",
		INIT_3D => x"11DF784E98E3A3133EB7B075B348235CACDC4DF712870F8AE111EC6169DF3673",
		INIT_3E => x"DD8BCD0DB05B4252F21FEE98ADBFB329BE08B7C5BD9891D4C8ECC8A80E8271A6",
		INIT_3F => x"11111111111111111111111111111111ADDF0BDF563CCA4C08AD132007D46503"
	)port map (
		DO   => doutout,			-- Port 16-bit Data Output
		DOP  => open,				-- Port 2-bit Parity Output
		ADDR => addrin,				-- Port 10-bit Address Input
		CLK  => clkin, 				-- Port Clock
		DI   => (others => '0'),	-- Port 16-bit Data Input
		DIP  => (others => '0'),	-- Port 2-bit parity Input
		EN   => '1',				-- Port RAM Enable Input
		SSR  => '0',				-- Port Synchronous Set/Reset Input
		WE   => '0'					-- Port Write Enable Input
	);
	-- End of FRAME0000_RAMB07 instantiation

end FRAME0000_B3;