--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
--	Grupo de Apoio ao Projeto de Hardware  - GAPH
--	Projeto X10GiGA - FINEP/PUCRS/TERACOM
--
--	M�dulo:	Mem�ria - Gerador de Frames - Prototipa��o
--	Autor:	Jeferson Camargo de Oliveira
--
-- 	FRAME:	0003
-- 	RAMB:	01
-- 	CONJ:	A
--
--	M�dulo gerado em 17 de July de 2008 �s 16h55min pelo
--	programa gerador de frames OTN do projeto X10GiGA.
--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

----Pragma translate_off
library unisim ;
use unisim.vcomponents.all ;
----Pragma translate_on

entity FRAME0003_A1 is
port(
		addr	: in  std_logic_vector(9 downto 0);	-- Barramento de endere�os da porta
		clk		: in  std_logic;					-- Entrada de clock para a porta
		dout	: out std_logic_vector(15 downto 0)	-- Sa�da de dados da porta
	);
end FRAME0003_A1;

architecture FRAME0003_A1 of FRAME0003_A1 is

	signal addrin	: std_logic_vector(9 downto 0);
	signal clkin	: std_logic;
	signal doutout	: std_logic_vector(15 downto 0);

	component RAMB16_S18 is
	generic(
		WRITE_MODE : string;
		INIT_00,INIT_01,INIT_02,INIT_03,INIT_04,INIT_05,INIT_06,INIT_07,
		INIT_08,INIT_09,INIT_0A,INIT_0B,INIT_0C,INIT_0D,INIT_0E,INIT_0F,
		INIT_10,INIT_11,INIT_12,INIT_13,INIT_14,INIT_15,INIT_16,INIT_17,
		INIT_18,INIT_19,INIT_1A,INIT_1B,INIT_1C,INIT_1D,INIT_1E,INIT_1F,
		INIT_20,INIT_21,INIT_22,INIT_23,INIT_24,INIT_25,INIT_26,INIT_27,
		INIT_28,INIT_29,INIT_2A,INIT_2B,INIT_2C,INIT_2D,INIT_2E,INIT_2F,
		INIT_30,INIT_31,INIT_32,INIT_33,INIT_34,INIT_35,INIT_36,INIT_37,
		INIT_38,INIT_39,INIT_3A,INIT_3B,INIT_3C,INIT_3D,INIT_3E,INIT_3F : bit_vector
	);
	port(
		DO   : out std_logic_vector(15 downto 0);	-- Port 16-bit Data Output
		DOP  : out std_logic_vector(1  downto 0);	-- Port 2-bit Parity Output
		ADDR : in  std_logic_vector(9  downto 0); 	-- Port 10-bit Address Input
		CLK  : in  std_logic;			 			-- Port Clock
		DI   : in  std_logic_vector(15 downto 0); 	-- Port 16-bit Data Input
		DIP  : in  std_logic_vector(1  downto 0); 	-- Port 2-bit parity Input
		EN   : in  std_logic;			 			-- Port RAM Enable Input
		SSR  : in  std_logic;			 			-- Port Synchronous Set/Reset Input
		WE   : in  std_logic			 			-- Port Write Enable Input
	);
	end component;

begin

	addrin <= addr;
	clkin  <= clk;
	dout   <= doutout;

	-- FRAME0003_RAMB01 instantiation
	FRAME0003_RAMB01 : RAMB16_S18
	generic map (

		-- The following generics are only necessary if you wish to change the default behavior.
		WRITE_MODE => "NO_CHANGE", 	-- WRITE_FIRST, READ_FIRST or NO_CHANGE

		-- The following generic INIT_xx declarations are only necessary
		-- if you wish to change the initial contents of the RAM to anything
		-- other than all zero's.
		INIT_00 => x"C027B9B7847C10C40BE3A13C17EB624E5F4EB3308A68EEA58C7AAF4005D2F628",
		INIT_01 => x"A1AC6400AA66F05C860E74E565FFFDD3943D5C59063F2ADCA8A00817AE9BD62F",
		INIT_02 => x"00EEB8227AF2586161E2EC50899D9610A86E6FACE660CCE0D8DDCA22FA4CD8B4",
		INIT_03 => x"C997F46836E1868D8BC2B526B933EFF8FC5668BF1F3DA1D88DB5700173CD6565",
		INIT_04 => x"0629F1EC5236B4898E0537B8864457DB567C038B9F1B5610E61E4C8633F28DC3",
		INIT_05 => x"1B4A29653C14E022D9E69DCB11CB1099E2D62BC02C944F2F365E14A78BFA9385",
		INIT_06 => x"0ED50BA3E5CCE17A4FCCABF09422C636BA3832AD1D0895DE373C98740C187774",
		INIT_07 => x"47D7661A5E9C4E2FAC36346ADDE50CDAAE580F7B32841D3595699A209149F199",
		INIT_08 => x"4B23D838F817BD2C7D8525D7F4ED52C64E310BFD82D944A07B1564DDCD823240",
		INIT_09 => x"D4C75A9D85EC4ADC4DE8E3B72489ED316007C518CDD17FF8EF71F1BD2A1A08F9",
		INIT_0A => x"041687064671E0EE074C60356AD57EDC5B8EFC5A0AAFF0B581565040B11A49DC",
		INIT_0B => x"26E919AE78BB934443F4A7CDD94119B75096FE6218689242E7A18FFF70D63227",
		INIT_0C => x"F812B002E5159CC483F7A55F746CE9A34E60FF7868A4A729B80B07440A642D89",
		INIT_0D => x"B051435FBC19ACC4486775F7301BB9402117E80E2318526611DEF57C59C33898",
		INIT_0E => x"4D9D553A6424FC92C90798EAF33981483F9E9ECDC0783489198A1649EB507EAF",
		INIT_0F => x"F8E6C4F66A5C5D233477E71DBE24EA2CC4AC6EE926161E72C144B5E0CDEEC355",
		INIT_10 => x"0AAEFFBDE7603602AC03D55B77B9F58B89B226E0177D04C50938FCD55615D2DB",
		INIT_11 => x"00B9F9DD2C70BB13D716F89DC96E165AB92C1504F26F3D8450D64D87969EE0D9",
		INIT_12 => x"A460A7E1A9DAC1BC58DDEF00F07AE6AAD0E6DD5BAEFDA01CFF861A876E592DC8",
		INIT_13 => x"FBEEDA8DC1FF00208E4F0D5CC00802F5C847785E738E60298B23CAD1FA449A9D",
		INIT_14 => x"599B748F607164C94D240AB6B10F8495C13CDBE8A75521C7A5BA9DA7263FBF28",
		INIT_15 => x"C5873588CF2759C76E6D5692670C1DBC014A2902E2C645792D762CB2E48E870C",
		INIT_16 => x"819AF5D74A0C249D6C9C68A84A4265DED6581F33D13252C077037EDAFD6B29F7",
		INIT_17 => x"97D7649B460CAB78D309122F435D4CA1164CC19FAF4251C454C9B4079DDD9328",
		INIT_18 => x"4FB07888E1542F132B8EE3863B2F249356915677D3AF7699B09D35C4DC8CBAC2",
		INIT_19 => x"A12CE930AF3631E7FBEFAD8CA3893A2D15B7BBBA0BC43185BF83C79E3CA93505",
		INIT_1A => x"8010DF3D6B74C5147CA72447054274615993946A5892A2C7AFD96CF712D78450",
		INIT_1B => x"3DDA81364B2C86346E707CB487AB28E9253E8015C46F73D5CC6B641240C705BB",
		INIT_1C => x"6615B9C7D3F7A56ED53DCE3228693960563618D501A2B57E818CD6945EA7E783",
		INIT_1D => x"90A1E9506FC51043CB8AA6F3503E35FC9E096CCF66EFC08657401BC2886BC488",
		INIT_1E => x"48AADA97C7905F4425CA0D6654A8B12C4A55E2FCC6138C29878CF6F2EAFF7850",
		INIT_1F => x"7452E9E633403594961DEBE9C605F43B961FA946E32ECB68CBBB929595664EA7",
		INIT_20 => x"D4A5FD928905A3C4DDDE0C4706C626450E3324715FB5BCA0EB8AEF0B1CE0A1A4",
		INIT_21 => x"8451EC85390044011C6DA9819F23B0E7BAA33E0DAC232BB288DD050F12321355",
		INIT_22 => x"FC6A83F058344ED76E6F613A0ADA4DA75F74E1B40E6EF4994B0D580A998CD77C",
		INIT_23 => x"DAD0281AAB43776ABCE92CAAA672AEA7573BA383A8499131C0B00E5111D53ABB",
		INIT_24 => x"A008886AA2928F2F15C94A67C54FC29EB5D56C9B8B5306B4B473EA0FA9E76E02",
		INIT_25 => x"4642AB746298174F1D2259894EDE87DB6D337582E218597479F99012601A6844",
		INIT_26 => x"C851673A6693A97E5DE02122B8B351DCA59E61F96DA79FBD32EA9E86D02E2245",
		INIT_27 => x"6C377BE7616A1528E77AF3FD97AE32BBD55ED846FFDFBFBDFF0A1C215F9827B1",
		INIT_28 => x"1605644555E07D26BACEB485E41F274D19F544AA49496AEB8AD3D6279BD190DA",
		INIT_29 => x"7E86914264DCC00A6BF262BC3FBBA4523BFBE1BB2F68AB130E29EBE174ABF28F",
		INIT_2A => x"C6745699DC92C77017C9A1F834463CCBACA7818D3FBACCFAF56A3D22B54B8863",
		INIT_2B => x"B333FE16CFAF2AC8F0631E99DEA40FD90A8A59C65AAC21848C56BDB2613ED575",
		INIT_2C => x"64D0DD4B5A341429A66341126BDD781B64A8938709CA34FF2D027737AC2C6E2E",
		INIT_2D => x"6E8AEF9FC452B5E2CC451C51C40BAD95F68D7F5FCC924DFC0F210BFBEA2D8DBC",
		INIT_2E => x"90DF9BD4D92023FD5A2495BB7EAA02760DB895DC2ADF197CE5F0C88D65AE21BA",
		INIT_2F => x"D76FE9B14462F0721E8EDD8CE3E1ACDC482271DDE5B8175280B9FE506EB880A4",
		INIT_30 => x"7C448978C1B8261AFFFABFEA5A7804FF89D89D7BDF3DDBA90EA4AB463ABDCB93",
		INIT_31 => x"A2355C69849769884035B01AAD9453469BD71A3F2DBF85DAA825CF4033C5CE30",
		INIT_32 => x"CF88D8956BEE18239EE0F39A3DE73494BFC4E04DA502180C5E14356A2982BF0F",
		INIT_33 => x"34C564EA82DB7CD3E3775F8EEAEC8D0322509FADD0D6D8401AF64899C8CD0288",
		INIT_34 => x"83A988B64105BED83D00EFACF7CC88CD1ABBADB60770639292C1BBD6F4E11FDB",
		INIT_35 => x"B038F30FE18BCCED18FC18EF3B1FED5012C37F5007CFBCB8A91E90C82C76EDB6",
		INIT_36 => x"7901918CC22EF76E6175F13EFB31FD13219E25E9BEC4BA035CA1AA3E55BB4231",
		INIT_37 => x"7488D7E5A1DAEB1755129356794AF44520A60348016E9C11E34BCF026AAB10A4",
		INIT_38 => x"B52068C149BBBC114491B4FA91A13500C1EECF98A46D5A1823B7359D64838AD6",
		INIT_39 => x"D19C6290115470C3ADF6CB84CC799A77E89628592509F594F2F56E0E30EA1D1E",
		INIT_3A => x"4D4E808CED5A9D41FA134E1CB12B43D9D8392217CB04269C182E8DE30ED0E213",
		INIT_3B => x"11FC9F578B39FF2DB06932DDA4221A5E1E64D462241D5B474A7DFA74A2131031",
		INIT_3C => x"071E8A76D04533B6B6779089A75FF8E9C5ADF40C049B63E58E37BDF8194EB50D",
		INIT_3D => x"CD26525AEDA5A49C881EFA2485874B60CED11649A16ED007A1A4B0DA18D477FF",
		INIT_3E => x"25129870F5488946C818CD20A52FFEDF222EBCDD7B64F51D1EF35FA369230035",
		INIT_3F => x"47E4088BCAF9B26D38A777922F3B104F93D74C7EB2CD63A0B3BA72A892D57881"
	)port map (
		DO   => doutout,			-- Port 16-bit Data Output
		DOP  => open,				-- Port 2-bit Parity Output
		ADDR => addrin,				-- Port 10-bit Address Input
		CLK  => clkin, 				-- Port Clock
		DI   => (others => '0'),	-- Port 16-bit Data Input
		DIP  => (others => '0'),	-- Port 2-bit parity Input
		EN   => '1',				-- Port RAM Enable Input
		SSR  => '0',				-- Port Synchronous Set/Reset Input
		WE   => '0'					-- Port Write Enable Input
	);
	-- End of FRAME0003_RAMB01 instantiation

end FRAME0003_A1;