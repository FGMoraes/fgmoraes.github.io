--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
--	Grupo de Apoio ao Projeto de Hardware  - GAPH
--	Projeto X10GiGA - FINEP/PUCRS/TERACOM
--
--	M�dulo:	Mem�ria - Gerador de Frames - Prototipa��o
--	Autor:	Jeferson Camargo de Oliveira
--
-- 	FRAME:	0003
-- 	RAMB:	03
-- 	CONJ:	B
--
--	M�dulo gerado em 17 de July de 2008 �s 16h55min pelo
--	programa gerador de frames OTN do projeto X10GiGA.
--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

----Pragma translate_off
library unisim ;
use unisim.vcomponents.all ;
----Pragma translate_on

entity FRAME0003_B3 is
port(
		addr	: in  std_logic_vector(9 downto 0);	-- Barramento de endere�os da porta
		clk		: in  std_logic;					-- Entrada de clock para a porta
		dout	: out std_logic_vector(15 downto 0)	-- Sa�da de dados da porta
	);
end FRAME0003_B3;

architecture FRAME0003_B3 of FRAME0003_B3 is

	signal addrin	: std_logic_vector(9 downto 0);
	signal clkin	: std_logic;
	signal doutout	: std_logic_vector(15 downto 0);

	component RAMB16_S18 is
	generic(
		WRITE_MODE : string;
		INIT_00,INIT_01,INIT_02,INIT_03,INIT_04,INIT_05,INIT_06,INIT_07,
		INIT_08,INIT_09,INIT_0A,INIT_0B,INIT_0C,INIT_0D,INIT_0E,INIT_0F,
		INIT_10,INIT_11,INIT_12,INIT_13,INIT_14,INIT_15,INIT_16,INIT_17,
		INIT_18,INIT_19,INIT_1A,INIT_1B,INIT_1C,INIT_1D,INIT_1E,INIT_1F,
		INIT_20,INIT_21,INIT_22,INIT_23,INIT_24,INIT_25,INIT_26,INIT_27,
		INIT_28,INIT_29,INIT_2A,INIT_2B,INIT_2C,INIT_2D,INIT_2E,INIT_2F,
		INIT_30,INIT_31,INIT_32,INIT_33,INIT_34,INIT_35,INIT_36,INIT_37,
		INIT_38,INIT_39,INIT_3A,INIT_3B,INIT_3C,INIT_3D,INIT_3E,INIT_3F : bit_vector
	);
	port(
		DO   : out std_logic_vector(15 downto 0);	-- Port 16-bit Data Output
		DOP  : out std_logic_vector(1  downto 0);	-- Port 2-bit Parity Output
		ADDR : in  std_logic_vector(9  downto 0); 	-- Port 10-bit Address Input
		CLK  : in  std_logic;			 			-- Port Clock
		DI   : in  std_logic_vector(15 downto 0); 	-- Port 16-bit Data Input
		DIP  : in  std_logic_vector(1  downto 0); 	-- Port 2-bit parity Input
		EN   : in  std_logic;			 			-- Port RAM Enable Input
		SSR  : in  std_logic;			 			-- Port Synchronous Set/Reset Input
		WE   : in  std_logic			 			-- Port Write Enable Input
	);
	end component;

begin

	addrin <= addr;
	clkin  <= clk;
	dout   <= doutout;

	-- FRAME0003_RAMB07 instantiation
	FRAME0003_RAMB07 : RAMB16_S18
	generic map (

		-- The following generics are only necessary if you wish to change the default behavior.
		WRITE_MODE => "NO_CHANGE", 	-- WRITE_FIRST, READ_FIRST or NO_CHANGE

		-- The following generic INIT_xx declarations are only necessary
		-- if you wish to change the initial contents of the RAM to anything
		-- other than all zero's.
		INIT_00 => x"30693F2AED8C74669AF86805B2A6A7469BD2A759A14B462377C84C51E93D9F33",
		INIT_01 => x"0B8467EA7D8072123A704D64F9DF21BADF0F45DACE4388891D4B82C8D7F33B72",
		INIT_02 => x"3A6300A150D0968AF96CDC79D704A063B54457ECDF123783379B67CD699DF558",
		INIT_03 => x"E7C3138E3A49EF6767114485B1385C16881E391BD527F561CF70414AFEF2648C",
		INIT_04 => x"6897953433DE081ADE0C6AAB36A8635A8F9E7FC71B0CA8B19875B5D11EF9D333",
		INIT_05 => x"25F3162E88470FFAFF7656073BE186B021A19DB6968B260E5DF013EB10A11A0E",
		INIT_06 => x"D184C8A540ED872EEF4558DC3CC4F3586D7700C7F99A7D78FC2A5BE18F3E97EA",
		INIT_07 => x"C4FCEA613C0BA29751FFFA1479D4EC6FE660CE95EEA5D59AAECFE847E52A3DCE",
		INIT_08 => x"16515902AAF0C7BCB1DE801BD7D7905D74180F141936F53E9081E93B60C980E7",
		INIT_09 => x"DB8553BE66050EDE86254372F50C903B826F2F3420755B42CC3CD3188DA1F9C9",
		INIT_0A => x"C3EB7B83D3AA683546AEF0090C3CE2D0D70C1A0C9BAB178450C60996C4110711",
		INIT_0B => x"7A2C8641C992BEDF249CAEC3B810A23ECF416C72BCF8703AC473A18FCE4436AE",
		INIT_0C => x"324049914E26B32F03F34DB949A1774B9190165B595B914AFFA5368F5E26258C",
		INIT_0D => x"20E2E53E9E82D980D701B1876199420DE2B84AF54DC53F578F55DD78FF68C611",
		INIT_0E => x"13B2B479F6A563B7ED6011B63872DB27B84C43282F296F004C7CCC4716AF22EB",
		INIT_0F => x"1499BDB44B9E3B1DCD67307E1FBF39FAC8C654F336EC1EF05A78CE581EA3240A",
		INIT_10 => x"2DCA491E1F9E5DEBAA8612563A8B0E8E5F35FE55CC474D0ECAF5BA673697B368",
		INIT_11 => x"C9D55557AF0189B8C9094FFDF216FF4A6182BECAC5CECCEDB9924987F838DF0F",
		INIT_12 => x"22322E4D320834C8399CAE81BD4F4986DF428DF3E24B5E3A3AA6B90B5B8D53D1",
		INIT_13 => x"A9E9B6D9B3770BDF09D640E1790E0039880BE61980B48B842DE522649A216BB7",
		INIT_14 => x"0F3CFC0C7DCAEA06E2DBFAAFDF941C5D8BD8CFEE8F1026BF011719D9BDE673ED",
		INIT_15 => x"93C06AB939A898A501658DB5F5F47F6199A799889DCD5D84B8DFAD761E2330CC",
		INIT_16 => x"74B1864B9AE7B5BEE66E51D748E3ADE060CEBFFAB441EF8D4A54CFB721F8F460",
		INIT_17 => x"392397ADD72FC0271C54349E7274432521FD30657D174ED78855E66BA7E6CEF7",
		INIT_18 => x"68FCA33CA96558C97A6C363A4BD8A14EF07241E808A582AF3A209B99CAE1C748",
		INIT_19 => x"B0DBED473D2B1A4228AF3A82FDD15432A1A9381604FEAE5BAF49E16A63DF29BB",
		INIT_1A => x"D2EBA43FA1CA8F8BB8B3512DA8C5759EAF84ECAFCC02CF8555A06919DC18A1B3",
		INIT_1B => x"398B26A41A30613C6F5CD71475A8B7C1D2A7C61ECE784CED5C07987CEF45DF72",
		INIT_1C => x"5F09A8E06A0C3697FEF65A3EAA7929B0B761C1CBFFBC8BAAA4C1AEB5F02C1E73",
		INIT_1D => x"40F58F8C32115EDD09056EC0E84F2039BA01E752E5E394AD5B7C4C21C1EF8C3E",
		INIT_1E => x"03E8D0418FB18820EBA600D4E3E89F98875B2868F0C06A0B6D2B32EB48027415",
		INIT_1F => x"8252DF189BF25925287C2A7D18B37D90BCA6B6EBA1A54159D3E6520555AB2941",
		INIT_20 => x"1BCF8B7224C4534419DB124E9C31E5285D250DF80EB9168047390323C9E46813",
		INIT_21 => x"AC2658874DAF8B2F75FB9D2015774FB30F90A9BEF37C7E4E054070747F85B12E",
		INIT_22 => x"3E52172D969DC599ED7C08DD0D08CFA62D5796262A69DCEF586C7FA7C444AA05",
		INIT_23 => x"DB23F96CEC7D50424F698D0F90EA3E080B1BE752D08625F46EE95A3C5B4F03F2",
		INIT_24 => x"B68BE1DC14305A7DB0E08D3F1F35011778539B594BEE2942DE7A0C4E55E543D2",
		INIT_25 => x"88C8F93C31B60A7B669F84D0226E66DFB555B85944DA9BD26ED508878F8A236B",
		INIT_26 => x"4DA3882E8103B34E65AA2BF5B3C1E42B358AF93D863EA8C6613ADC0B4A48A617",
		INIT_27 => x"442D6B546B02C4204642A7F44315CC3E1D20FC7EE32B60D2B453C6B550B54A4F",
		INIT_28 => x"88EC8877941645705F84DD7FD66B552031E498E36FBD9CBED9111A2D80D446CE",
		INIT_29 => x"8C9BDA24080E8E43811B19002C065FCC04E0CBD798BC6EC384D6D31DF61E1DF5",
		INIT_2A => x"FAB916EEE4E195CEF19663ED80373A5244C02753C5D6E2D3CE58C49E91B5F593",
		INIT_2B => x"28B0A131F2F4D8FA1E542A196110D3048108C9033DEA46F322F2D6F5F0406B0D",
		INIT_2C => x"83342BF670D04245477CDB831E865D0B165F2FBDEA1A3A46C9404266318994DD",
		INIT_2D => x"1F841672ADA61F575F1B0F9235AA7320AF44ABFD732D2BE4583388446757C64D",
		INIT_2E => x"95F632703932F5930DFB66052FCB16BC4EA51CD7B3F5040D4EACA62BB31D6905",
		INIT_2F => x"1896644605ACB1CB05903BE7DE7496C95745CB4832482E84418AF76C3A1623CF",
		INIT_30 => x"E0EDD6624A5BCC74A7571A8A59C5F6FDA8F2125EBFF39D69E80DDF5D9DC4E960",
		INIT_31 => x"BE4708A7B6905A704D594AC69A0371CD6EF17B5E6EEA1C7B8A707E0750DBBE8B",
		INIT_32 => x"FBAA98F43FD9852C968471A9FDD6B0C1D72A9012803E01B99C8A56BC7B4128B7",
		INIT_33 => x"847008BF2333BEA3205BB2563F88F046CF682C9807D3735FFC9520FF61C9225A",
		INIT_34 => x"21FEBB89A97443DD13AAD1F8B1B69F0525F46872B812CDA9C2F15AA50D05753D",
		INIT_35 => x"07431368C927BB825A997999C75246EA889433D3F849A8520B43C4751D618FD4",
		INIT_36 => x"7753B03C7C1EF62CCB08A95CE042BB2138F28A02EEA88C2631634DF980AC7834",
		INIT_37 => x"A558904060382CCAD020727828D98C2BBAEA8129ADC0360E5F9548A6D2BEC6D7",
		INIT_38 => x"A2A84BEF2CA05F677BC6E1692F508E677AF8039F59794E72D215757A7A2094C3",
		INIT_39 => x"FE3171070A2B61F035EF3E037F5089480A707063F5230FE211EC43F84977F0C5",
		INIT_3A => x"771549D12E4D225AFAED43D4B24D9052D1FE534FB596764A83E6299C97CA2909",
		INIT_3B => x"E0509C286D9EB8602D97985C368E5A464A82BFF1CAA24280B447DBED11D7A4B0",
		INIT_3C => x"CD48E7ED0D4ABDF09A9B37B11A4BC382182AB29FC2D060543B0A22285FC3C53F",
		INIT_3D => x"BCFF5ABB1B15C9BA63A96DDCDA0981DBD0A9E1D1C8BBF5C80EDA912F6E61857F",
		INIT_3E => x"B684AF3ADCCDCB59D1B016B6CF9A42781C7AB44248E429D27B052B969DD8E066",
		INIT_3F => x"1111111111111111111111111111111130D257F05A83D2E89D5EEA2A9F5903F5"
	)port map (
		DO   => doutout,			-- Port 16-bit Data Output
		DOP  => open,				-- Port 2-bit Parity Output
		ADDR => addrin,				-- Port 10-bit Address Input
		CLK  => clkin, 				-- Port Clock
		DI   => (others => '0'),	-- Port 16-bit Data Input
		DIP  => (others => '0'),	-- Port 2-bit parity Input
		EN   => '1',				-- Port RAM Enable Input
		SSR  => '0',				-- Port Synchronous Set/Reset Input
		WE   => '0'					-- Port Write Enable Input
	);
	-- End of FRAME0003_RAMB07 instantiation

end FRAME0003_B3;