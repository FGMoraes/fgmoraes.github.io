--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
--	Grupo de Apoio ao Projeto de Hardware  - GAPH
--	Projeto X10GiGA - FINEP/PUCRS/TERACOM
--
--	M�dulo:	Mem�ria - Gerador de Frames - Prototipa��o
--	Autor:	Jeferson Camargo de Oliveira
--
-- 	FRAME:	0002
-- 	RAMB:	00
-- 	CONJ:	A
--
--	M�dulo gerado em 17 de July de 2008 �s 16h55min pelo
--	programa gerador de frames OTN do projeto X10GiGA.
--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

----Pragma translate_off
library unisim ;
use unisim.vcomponents.all ;
----Pragma translate_on

entity FRAME0002_A0 is
port(
		addr	: in  std_logic_vector(9 downto 0);	-- Barramento de endere�os da porta
		clk		: in  std_logic;					-- Entrada de clock para a porta
		dout	: out std_logic_vector(15 downto 0)	-- Sa�da de dados da porta
	);
end FRAME0002_A0;

architecture FRAME0002_A0 of FRAME0002_A0 is

	signal addrin	: std_logic_vector(9 downto 0);
	signal clkin	: std_logic;
	signal doutout	: std_logic_vector(15 downto 0);

	component RAMB16_S18 is
	generic(
		WRITE_MODE : string;
		INIT_00,INIT_01,INIT_02,INIT_03,INIT_04,INIT_05,INIT_06,INIT_07,
		INIT_08,INIT_09,INIT_0A,INIT_0B,INIT_0C,INIT_0D,INIT_0E,INIT_0F,
		INIT_10,INIT_11,INIT_12,INIT_13,INIT_14,INIT_15,INIT_16,INIT_17,
		INIT_18,INIT_19,INIT_1A,INIT_1B,INIT_1C,INIT_1D,INIT_1E,INIT_1F,
		INIT_20,INIT_21,INIT_22,INIT_23,INIT_24,INIT_25,INIT_26,INIT_27,
		INIT_28,INIT_29,INIT_2A,INIT_2B,INIT_2C,INIT_2D,INIT_2E,INIT_2F,
		INIT_30,INIT_31,INIT_32,INIT_33,INIT_34,INIT_35,INIT_36,INIT_37,
		INIT_38,INIT_39,INIT_3A,INIT_3B,INIT_3C,INIT_3D,INIT_3E,INIT_3F : bit_vector
	);
	port(
		DO   : out std_logic_vector(15 downto 0);	-- Port 16-bit Data Output
		DOP  : out std_logic_vector(1  downto 0);	-- Port 2-bit Parity Output
		ADDR : in  std_logic_vector(9  downto 0); 	-- Port 10-bit Address Input
		CLK  : in  std_logic;			 			-- Port Clock
		DI   : in  std_logic_vector(15 downto 0); 	-- Port 16-bit Data Input
		DIP  : in  std_logic_vector(1  downto 0); 	-- Port 2-bit parity Input
		EN   : in  std_logic;			 			-- Port RAM Enable Input
		SSR  : in  std_logic;			 			-- Port Synchronous Set/Reset Input
		WE   : in  std_logic			 			-- Port Write Enable Input
	);
	end component;

begin

	addrin <= addr;
	clkin  <= clk;
	dout   <= doutout;

	-- FRAME0002_RAMB00 instantiation
	FRAME0002_RAMB00 : RAMB16_S18
	generic map (

		-- The following generics are only necessary if you wish to change the default behavior.
		WRITE_MODE => "NO_CHANGE", 	-- WRITE_FIRST, READ_FIRST or NO_CHANGE

		-- The following generic INIT_xx declarations are only necessary
		-- if you wish to change the initial contents of the RAM to anything
		-- other than all zero's.
		INIT_00 => x"92E18271910C9089B49AE5FF33CE5F7D7FD28CE2653F5B641F861A8D4E91F6F6",
		INIT_01 => x"A2DF541B4703BA12056BAD202A5D6A311D31112ED8EC86398089A3C66BED0FBF",
		INIT_02 => x"7015519B8BFD91344D968CC019AFE26B7736DCBBEFCDFF905D07C1B303FA9D7E",
		INIT_03 => x"F093FD193CD2024368760E26DEF17D57D34E7826C6BCB65D02AD553474DF8343",
		INIT_04 => x"E797453372A3E88CC206855CD9B67268410DAC14F1FBE2CCAB52D971C4555D3A",
		INIT_05 => x"7721E15A041EAA326DC89C21940D5FDAC4D230D00367EEA73445701A4C7DEDBE",
		INIT_06 => x"0D1B5863FA60B1E1CC509A91F8ECD35404A0FEF7E4DAD2001C5E38937471B1AF",
		INIT_07 => x"805E8565B8716CF8976C9C06D2BA5454312D2141AF8BF5E4064E95CA112E8ACD",
		INIT_08 => x"65606EE0F94ED61263A8C5C49E8D45693A6FD7F24A6960930448A0F9F4420DE0",
		INIT_09 => x"DF02B21A410E64E5B66B3B157196208273A1B2319913E3F6EDEB49D32EC7990B",
		INIT_0A => x"0835D8966A66C7A597B25003990BE78BDB8866C486D29CF5B86599779F5F2AA7",
		INIT_0B => x"3409285895F782C9D0F362B81817E4EDA21B431E175FC4178DC08A60CF566667",
		INIT_0C => x"33B6B28C85D8761B1282B2532359B0DB84DFB0C66D44FB93DF90FDB33A878190",
		INIT_0D => x"6D67569F4C06FEAE18A0C4AFB301881B4D4BF4441EAE810A89FBF90D858167E8",
		INIT_0E => x"98E954C60C2C0D39347A85C51500209468E534A97551BE5B3D19FCE65E52A243",
		INIT_0F => x"DF39065AF0AE0142C0D7899A17C27296D1FAC634482F9E727904AFA8A2798100",
		INIT_10 => x"E85CDB04EAC585F376BAF4586E13082FC0269E444D542913D1E06E4251D484EB",
		INIT_11 => x"D78878DB5C4775CF90A5087B8D47A859CAB974CBCDDA6C90F77BFE5CA56BBD7C",
		INIT_12 => x"C52C7403249B508EA88928225ABB46767230F374099A4A9706F665D2A7C16B4C",
		INIT_13 => x"6461E883561A52EC28BEC151797262038B9F21A7E81F4EDE7386EEF181C4BFA3",
		INIT_14 => x"12CC20DD90F8B807476CA194666F223B0289BEFC0289C765F7AA480EEC7473B4",
		INIT_15 => x"17CD5E2DEC98DB7E0DC23384501481AF06048A8C5A2546836A64BF4865F14345",
		INIT_16 => x"5E3DCF6351AF6D042535BF3D5F641C21FC6EDB50E92EA6F483B65483F6E25DFF",
		INIT_17 => x"32F30E0E4014BB87BE42D9322EB2C0DBEB1E39A6FA3198F1CCFEDAF3030C09F6",
		INIT_18 => x"4B7D2F848897017BE48224C646574EA590825ABD07CFE5DB29A0ABBE49F834AF",
		INIT_19 => x"FBB84839EA35B65246D66BDEAA07ADE3E1EEEFC7C26E19CDD2F789968827C6BC",
		INIT_1A => x"40E2367ADE6273159AD8D5317066E631235E29B65B38F521333F29554F31082B",
		INIT_1B => x"E91D425C19295EA17934260A29DFB91811718C3A52AD779E8DE14A6D8680BAE5",
		INIT_1C => x"FF8162650BA4A769612EB2426169492580D58C98596C8A769E40E65D6646445B",
		INIT_1D => x"57D73DAD9F3FAC3610DB67630DF4362E122C2B0EEAEDB8D0CA2A4AC7FF9FCB9E",
		INIT_1E => x"33A979045CAA359D88D2B38EE3033B25D1C0DDA5662356F34388D8C3E33EDC56",
		INIT_1F => x"E3C3B557070E42B5267E4D2F42BE019139D2EBBE075B20957DD52B7D09928897",
		INIT_20 => x"1E72530CA4D8FC6D050ADBE9707AEBA8C801B4609CB3C2A59F412B7826D2B568",
		INIT_21 => x"259159BFF7FEDFC569601922E466A138032F21E87986F510C2ED2D72469E1E67",
		INIT_22 => x"4068EBCCE3FC07F1CE86D9A1D56483F424EB3ECA9447ED72B8B1DB5E9CD2B1BC",
		INIT_23 => x"C7661751BC4E04E8C56A78780F6387624042D4EC6D6C4EC785191F35EF8EB0B9",
		INIT_24 => x"E2F7649F9C969F52E1EAB0B7E35D1488405EE9C3B6237516E70C29D8E5E0D3EB",
		INIT_25 => x"706164C23099EC1D4B7DD8A31027046308820257AE9C8DAE740B52F7D0F30758",
		INIT_26 => x"6E075573AE42FC5B2E5E6CA17D59FB15E3CB30466150BB6931C323CD3D1EEA6E",
		INIT_27 => x"77B3B8DE2010C3FB1DE5B59CD1F6E5F292DE74D9B8C6F8353FC1F77EC6235E47",
		INIT_28 => x"1C99B49744964CD12654E6C03E75F28C93A18748B71B8E04D12585D46453ACC3",
		INIT_29 => x"52E263AF69BAAD837341A41BD6124356363BD9FE9DF90EC74ECEF0BD4F57066E",
		INIT_2A => x"DC98DC564EBAE73323FB96DFC8A418505001953270F8590AD0490171C929D4D6",
		INIT_2B => x"886BB02516E3FFAA988B33164ABEB9D1B3B06C6B9F1FC616B985DF2844C9E35A",
		INIT_2C => x"E1D01FEA7033F40B3B05F9CFD6B988F4DA067743E3737A63A5DB17AE702B3FF0",
		INIT_2D => x"B71DAFCBA866D787157A627DE0EA8BA01025E79BA7EF1510872CCC974F933769",
		INIT_2E => x"3E2A1767D4306BE23B69D9F30FB6DFC92D6DE4935D48F3BCCD3878F984FC45EC",
		INIT_2F => x"DBEECD52ADDDFFE7918AABD77C51D3B87DB0DFE834A6B2E813AB71EDBB3E2848",
		INIT_30 => x"3EB30BC9A20CA4B748332278152E063FA8A1D0B787455E0BBAE712A0749EDDDD",
		INIT_31 => x"4AA3E4704DAC6F7E6748C7106684BAEBB69A02FD4C1BB4D9EB2173A7F1FC31FB",
		INIT_32 => x"0A6DC809B16F308C4FEB5E2C77823983F0D47C8738414BB0B79564C1E086E52D",
		INIT_33 => x"A02DC7460F79E5394BBA1928B47D6ABCF0A3D748D86D34D11920A7AE79625A23",
		INIT_34 => x"A3E00D4DBED9093F9BD810DAF88B53D571B2281832948C9B930DFE8B5B511C1E",
		INIT_35 => x"1BAF93D86A271C58D48597DAB402302AF806A5C8A3CE6B0EE9CBBEDBDB249EDB",
		INIT_36 => x"9EC2023689735AC2AF59E17E8B2518CA4DFCA8BB3E93C6E1817F92A318B1A977",
		INIT_37 => x"D83ACFA09DD1661977F4DDB52033AA5D05CF5F37877954DCE3CB43A95C1D7AE2",
		INIT_38 => x"3BC7770852BCCE42E3A6D212AF97AB378A0B96B38464667526513770EED2FB75",
		INIT_39 => x"FE8A846DB48BBF904BF8D1143CD8C8ACD7A616855914CF180C3AEF026831892C",
		INIT_3A => x"2E1B7A7D892A41B80B578CD9D80712A4DCFCE00BA4ED04E165F14996E896D213",
		INIT_3B => x"B02FC30401FAD9A7BB6A4691668C5CDBC72DF6564F1373F43CEFD7D4D7F045F8",
		INIT_3C => x"10073C7C83C1DA0A5A988E144D04E1CEC2D78A74685965C15AF0F693A911E09E",
		INIT_3D => x"703B47B59BE4F74BA6719B0B69B545C85E6F8B3D4C86A1BBF6C06B86D5287E22",
		INIT_3E => x"74D39DBF6721D28F4E84126AF7DBBE26066F481D28D848A82C2DF354569260AE",
		INIT_3F => x"38A6E36CADB6714256585526DFC1DDE344343A9CEFB1159A508304E9D7BB227D"
	)port map (
		DO   => doutout,			-- Port 16-bit Data Output
		DOP  => open,				-- Port 2-bit Parity Output
		ADDR => addrin,				-- Port 10-bit Address Input
		CLK  => clkin, 				-- Port Clock
		DI   => (others => '0'),	-- Port 16-bit Data Input
		DIP  => (others => '0'),	-- Port 2-bit parity Input
		EN   => '1',				-- Port RAM Enable Input
		SSR  => '0',				-- Port Synchronous Set/Reset Input
		WE   => '0'					-- Port Write Enable Input
	);
	-- End of FRAME0002_RAMB00 instantiation

end FRAME0002_A0;