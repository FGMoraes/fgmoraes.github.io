--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
--	Grupo de Apoio ao Projeto de Hardware  - GAPH
--	Projeto X10GiGA - FINEP/PUCRS/TERACOM
--
--	M�dulo:	Mem�ria - Gerador de Frames - Prototipa��o
--	Autor:	Jeferson Camargo de Oliveira
--
-- 	FRAME:	0003
-- 	RAMB:	01
-- 	CONJ:	B
--
--	M�dulo gerado em 17 de July de 2008 �s 16h55min pelo
--	programa gerador de frames OTN do projeto X10GiGA.
--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

----Pragma translate_off
library unisim ;
use unisim.vcomponents.all ;
----Pragma translate_on

entity FRAME0003_B1 is
port(
		addr	: in  std_logic_vector(9 downto 0);	-- Barramento de endere�os da porta
		clk		: in  std_logic;					-- Entrada de clock para a porta
		dout	: out std_logic_vector(15 downto 0)	-- Sa�da de dados da porta
	);
end FRAME0003_B1;

architecture FRAME0003_B1 of FRAME0003_B1 is

	signal addrin	: std_logic_vector(9 downto 0);
	signal clkin	: std_logic;
	signal doutout	: std_logic_vector(15 downto 0);

	component RAMB16_S18 is
	generic(
		WRITE_MODE : string;
		INIT_00,INIT_01,INIT_02,INIT_03,INIT_04,INIT_05,INIT_06,INIT_07,
		INIT_08,INIT_09,INIT_0A,INIT_0B,INIT_0C,INIT_0D,INIT_0E,INIT_0F,
		INIT_10,INIT_11,INIT_12,INIT_13,INIT_14,INIT_15,INIT_16,INIT_17,
		INIT_18,INIT_19,INIT_1A,INIT_1B,INIT_1C,INIT_1D,INIT_1E,INIT_1F,
		INIT_20,INIT_21,INIT_22,INIT_23,INIT_24,INIT_25,INIT_26,INIT_27,
		INIT_28,INIT_29,INIT_2A,INIT_2B,INIT_2C,INIT_2D,INIT_2E,INIT_2F,
		INIT_30,INIT_31,INIT_32,INIT_33,INIT_34,INIT_35,INIT_36,INIT_37,
		INIT_38,INIT_39,INIT_3A,INIT_3B,INIT_3C,INIT_3D,INIT_3E,INIT_3F : bit_vector
	);
	port(
		DO   : out std_logic_vector(15 downto 0);	-- Port 16-bit Data Output
		DOP  : out std_logic_vector(1  downto 0);	-- Port 2-bit Parity Output
		ADDR : in  std_logic_vector(9  downto 0); 	-- Port 10-bit Address Input
		CLK  : in  std_logic;			 			-- Port Clock
		DI   : in  std_logic_vector(15 downto 0); 	-- Port 16-bit Data Input
		DIP  : in  std_logic_vector(1  downto 0); 	-- Port 2-bit parity Input
		EN   : in  std_logic;			 			-- Port RAM Enable Input
		SSR  : in  std_logic;			 			-- Port Synchronous Set/Reset Input
		WE   : in  std_logic			 			-- Port Write Enable Input
	);
	end component;

begin

	addrin <= addr;
	clkin  <= clk;
	dout   <= doutout;

	-- FRAME0003_RAMB05 instantiation
	FRAME0003_RAMB05 : RAMB16_S18
	generic map (

		-- The following generics are only necessary if you wish to change the default behavior.
		WRITE_MODE => "NO_CHANGE", 	-- WRITE_FIRST, READ_FIRST or NO_CHANGE

		-- The following generic INIT_xx declarations are only necessary
		-- if you wish to change the initial contents of the RAM to anything
		-- other than all zero's.
		INIT_00 => x"968E1536AEC29ED6B7541ED287BC025C44D7A7E66D150A584B3116CB1CD6996E",
		INIT_01 => x"BE7A9BE88AC7A1C4B2EFF43D214B220A378EFB93E167DCD461757EC7B49FF0C5",
		INIT_02 => x"568F34F0FE01401D08941038010DACA75537094751B99BE48CF3BDBF05CB139A",
		INIT_03 => x"9DEED27BAFAC17E4E070D148357F9D358F2804F81E6FB9C6AA835BED7711640B",
		INIT_04 => x"6ECFB463F7E7589D74ECB0FE7EF27CCD09F2FB17A3BE83AE24F9C4542C330901",
		INIT_05 => x"9BD7EE6D3CBEBA85D64DD0112D6CA7A824F8D4916E9CDE64E4F9AB7579F27BCE",
		INIT_06 => x"5D11D2AA37AD98BA9CFE82C2D1C95500C7485401360F736B300478F57E0CB749",
		INIT_07 => x"C67971130357517BDEE2158CE24125105F8D617814E6E15A810B0E5801D45288",
		INIT_08 => x"8AC6FC113369DAE7F9AD25A5B8588324A9364B2347B4350040CA646F9D9AE6B8",
		INIT_09 => x"A4052FA56539505768C908A1657F4A55C7FE3F9CBC1E497DF53849B8149241CA",
		INIT_0A => x"0AD49A9E487C9FD0ED182794463E028D4F969D55ECAF4F432F0D39F2BB8A6676",
		INIT_0B => x"75C5DF832335468208644909CE37FBFEE9BDFCE7285C1123996E4EA22C8E3A47",
		INIT_0C => x"808458A9712B6F344A34104699C3048807631DDFAE6461AB104FCC18EBFED6E7",
		INIT_0D => x"B02C2B43DDA801DB25422A9F1FA8D5B9A9AF138BF479050B645D67597F08F3ED",
		INIT_0E => x"51A3CF3F221828E01B48F99998DFE47C37D1E1A39DC92C1525336533FB641E44",
		INIT_0F => x"46D1FBF8ADDAF6C05D2382417E74680F9F3F3CE602DCE03931861D17F731135E",
		INIT_10 => x"0CDF353A11762AB30BE4919FB698C11589167CDEBA498892A1B288E329C1323F",
		INIT_11 => x"E7A1ACBFBEC718131BF8633F35761A29816AD7CE783A7E34B35F23CB0263B4F6",
		INIT_12 => x"82A8DA6CD631D503287C86E019F3AF1F05A4191F9AEC58A6D65869CEC605933C",
		INIT_13 => x"45FE3CE15E342729B836CE3C5EB96E4DE2E95AEEB811A583847813B561A627E8",
		INIT_14 => x"7F9CFEC9B5C6DF0E3F273BBFE94C0EE6EE8CDEA5CB7F84C9A86009E49551D32C",
		INIT_15 => x"E71023F62C36277FB5F78BE03347A7D3EEED6F0EAA97B604CBFA4284588DC1A4",
		INIT_16 => x"D4171B7C140FC5A1ED3E019F95A5DCD831EA5ECCDE7C3EE29638D7B3B2BAC3D1",
		INIT_17 => x"10857BD60399E856E86F757C0C1DC963553CBC1066D0FF180FEC25805603AE9B",
		INIT_18 => x"23F8EC212986BDD9F1EA84013E32A4CEDC0CF3951D27D71AEE2FDECA1EA9B714",
		INIT_19 => x"600499BBB73B4862A3FDFD24BAFBBFAE874BED010FA59D6AF9D7EB9671FE80AE",
		INIT_1A => x"A55317DB80499A390660F24F6623FAF166F4DB9C36D844BC5AEA5AA53BF3D3B2",
		INIT_1B => x"4EDDA10B86D0E0350DC97C20A7EC43209640DE1B80D58B9AB9A07FE63B78632B",
		INIT_1C => x"A431EA80B0A10ECAE25E165EADFD180FF219AFB818042504D54374E2090B417B",
		INIT_1D => x"ED2E55255981DF08F6BB4DDD9F04CC30F9A9A5DB4359AF411FD371D99206B9C2",
		INIT_1E => x"8C8731E18AC7A9F03DFB599988B8EE38860CC49C4F769C692AC8C17D92C11601",
		INIT_1F => x"3C19E518601352EDAEB0E7FFE880A548495718DB31E4BC7882CFB433F7718F1C",
		INIT_20 => x"A45671DB2C579BC66EA93DCAC5F876B24D72540A75F82151D6C9756D3FC620E9",
		INIT_21 => x"9EB2B882A3BAE9C0CBAFE521C5AE5EBF05A4BD2CBD1A59911B548AC8E6E54B2F",
		INIT_22 => x"36755F848D2B131CBE4382C468D98C3CAF7AFC5B3E6B101F91F1A56821931D2A",
		INIT_23 => x"63E2470110102F8862899EFE2DFC759B3EA69EF26FD6608E660A5C324A273CB6",
		INIT_24 => x"9C4CDD1E310C47B64D6E9B0C22B462803D1713EB3304829C30BFAF4BAF1CECF3",
		INIT_25 => x"46EC750D536BD06C3F2D275C6D9D0B3D8B8B4DD7139E91632143235EF7CA04A6",
		INIT_26 => x"997B84F2C98683890E3A1ADA28736E74824C758898B411D6493E5EF00CD267CC",
		INIT_27 => x"652876192917B4489DCCB1EA7FCA9CEF70DF382EF5FF19EE1E6C1BD4409809D8",
		INIT_28 => x"866F2580B80CC34400D5A8D4A59CE3271EE0C2E6A2F1E1C26A72C6A9426A9DDE",
		INIT_29 => x"A42B224403016F2280A8F61EA8F2BB0554B7B90477D150AF49B29D73C55EE1FA",
		INIT_2A => x"8C8B7D091EF44D95CF00A6BA24CA9437BABEE74B80E21514C6BF629DE041A35B",
		INIT_2B => x"834F85FC15A900DAC32635F30888207AB7EA1A67F028C2E8D96DE64800AB982B",
		INIT_2C => x"8F901D2BF3E8ED73D0977E1198D6EA8DB8181EB432F3CCC0C09EC7FD3AF9CBCA",
		INIT_2D => x"EB19C72B52E5C491578C940BF9FB4DBD9DD8AA77BA53292147D650861CA65DFB",
		INIT_2E => x"F9E0AA9CAD27FBFCAAE0802719F1F67129FE7EF9B04C16FCB3A82A29BDEE67D7",
		INIT_2F => x"C9A98696AC7DB8B658F4A258C2439C9DAE3884DB42E239D7BC944ED3492422A7",
		INIT_30 => x"5F43E1203595CABF898D4F19D4B99CDD4B55420590E73782A87AB45C5AF34A4B",
		INIT_31 => x"4F7D77DD8CC384CA48A2F59252F430CF2C4CD87D6367F141A460197BB00E62D5",
		INIT_32 => x"B7429B72A8698D478B4039DFE4DD0A4E894A180A7DC0C35BD5DD61B75A100B49",
		INIT_33 => x"15DBB1FAAB8E2AEC6B6DDE3548FD11D1A69A49FDEE65FA41D8C28CE161E6FAEE",
		INIT_34 => x"38F92B76D079F923F40B5464BA7C6221CAABEFA227E4481BFFEE12DD9E700938",
		INIT_35 => x"85032D0892944457074EBB68841DFBB3CF984F2B0143CBB62B5BFE1DBFE2605C",
		INIT_36 => x"463DC7412117E282A5A530209D0CAB6D2B0E7B661E10773E8153DB000B315D12",
		INIT_37 => x"FB66FE304CB51441589F7AAF280D071271C224F78925B49CDA077FC9A00F2161",
		INIT_38 => x"94DBC384EE480D47CBB3638429108BFAC1B6C901DEB3DD337861725F1DD94EDE",
		INIT_39 => x"B97A7D45D80E60ECB204A6DB45646F865D59A44398A3EDB28EA4A3E93C7B67DB",
		INIT_3A => x"5C1E30B8CB4A8931EABA706ABC2625FEE482DC284DBE90F13743D28D545BEA78",
		INIT_3B => x"CA4DA1098F0C43B9BE588615882394A921D645AB52614F4DE3D0A26C314A1AF5",
		INIT_3C => x"ADB5E15D976C83A5A2F13FF5FF2B3EE43000CD1AEFB227420FCAC289ADAE5794",
		INIT_3D => x"C6DB28AA8F3102CA211667E1D7D26E6F2E51E203C00ABCAEF5A93CD69470B588",
		INIT_3E => x"9E3C7EF16E334D9F3281783F5EE7E1C2F49C51FD32D0DD6E133411F81BA9B60C",
		INIT_3F => x"111111111111111111111111111111117BEDB82D7D8CCF27085A08C9CAD520D7"
	)port map (
		DO   => doutout,			-- Port 16-bit Data Output
		DOP  => open,				-- Port 2-bit Parity Output
		ADDR => addrin,				-- Port 10-bit Address Input
		CLK  => clkin, 				-- Port Clock
		DI   => (others => '0'),	-- Port 16-bit Data Input
		DIP  => (others => '0'),	-- Port 2-bit parity Input
		EN   => '1',				-- Port RAM Enable Input
		SSR  => '0',				-- Port Synchronous Set/Reset Input
		WE   => '0'					-- Port Write Enable Input
	);
	-- End of FRAME0003_RAMB05 instantiation

end FRAME0003_B1;