--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
--	Grupo de Apoio ao Projeto de Hardware  - GAPH
--	Projeto X10GiGA - FINEP/PUCRS/TERACOM
--
--	M�dulo:	Mem�ria - Gerador de Frames - Prototipa��o
--	Autor:	Jeferson Camargo de Oliveira
--
-- 	FRAME:	0002
-- 	RAMB:	03
-- 	CONJ:	B
--
--	M�dulo gerado em 17 de July de 2008 �s 16h55min pelo
--	programa gerador de frames OTN do projeto X10GiGA.
--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

----Pragma translate_off
library unisim ;
use unisim.vcomponents.all ;
----Pragma translate_on

entity FRAME0002_B3 is
port(
		addr	: in  std_logic_vector(9 downto 0);	-- Barramento de endere�os da porta
		clk		: in  std_logic;					-- Entrada de clock para a porta
		dout	: out std_logic_vector(15 downto 0)	-- Sa�da de dados da porta
	);
end FRAME0002_B3;

architecture FRAME0002_B3 of FRAME0002_B3 is

	signal addrin	: std_logic_vector(9 downto 0);
	signal clkin	: std_logic;
	signal doutout	: std_logic_vector(15 downto 0);

	component RAMB16_S18 is
	generic(
		WRITE_MODE : string;
		INIT_00,INIT_01,INIT_02,INIT_03,INIT_04,INIT_05,INIT_06,INIT_07,
		INIT_08,INIT_09,INIT_0A,INIT_0B,INIT_0C,INIT_0D,INIT_0E,INIT_0F,
		INIT_10,INIT_11,INIT_12,INIT_13,INIT_14,INIT_15,INIT_16,INIT_17,
		INIT_18,INIT_19,INIT_1A,INIT_1B,INIT_1C,INIT_1D,INIT_1E,INIT_1F,
		INIT_20,INIT_21,INIT_22,INIT_23,INIT_24,INIT_25,INIT_26,INIT_27,
		INIT_28,INIT_29,INIT_2A,INIT_2B,INIT_2C,INIT_2D,INIT_2E,INIT_2F,
		INIT_30,INIT_31,INIT_32,INIT_33,INIT_34,INIT_35,INIT_36,INIT_37,
		INIT_38,INIT_39,INIT_3A,INIT_3B,INIT_3C,INIT_3D,INIT_3E,INIT_3F : bit_vector
	);
	port(
		DO   : out std_logic_vector(15 downto 0);	-- Port 16-bit Data Output
		DOP  : out std_logic_vector(1  downto 0);	-- Port 2-bit Parity Output
		ADDR : in  std_logic_vector(9  downto 0); 	-- Port 10-bit Address Input
		CLK  : in  std_logic;			 			-- Port Clock
		DI   : in  std_logic_vector(15 downto 0); 	-- Port 16-bit Data Input
		DIP  : in  std_logic_vector(1  downto 0); 	-- Port 2-bit parity Input
		EN   : in  std_logic;			 			-- Port RAM Enable Input
		SSR  : in  std_logic;			 			-- Port Synchronous Set/Reset Input
		WE   : in  std_logic			 			-- Port Write Enable Input
	);
	end component;

begin

	addrin <= addr;
	clkin  <= clk;
	dout   <= doutout;

	-- FRAME0002_RAMB07 instantiation
	FRAME0002_RAMB07 : RAMB16_S18
	generic map (

		-- The following generics are only necessary if you wish to change the default behavior.
		WRITE_MODE => "NO_CHANGE", 	-- WRITE_FIRST, READ_FIRST or NO_CHANGE

		-- The following generic INIT_xx declarations are only necessary
		-- if you wish to change the initial contents of the RAM to anything
		-- other than all zero's.
		INIT_00 => x"278CBC0EA9A5A66F97B16ABEA1D87197634C71E5CE93D5416970EB43D7672D83",
		INIT_01 => x"6F02503315DE79133268148105A647A1FDA5F6709993E9ACFEC5F4B8E6EA9028",
		INIT_02 => x"0B91C9541DFCF35F448971FEB0F199EF0448CF9A11A5B54FD4A00BCE7E39A513",
		INIT_03 => x"FA8A1D3CC9E17EAB8433859FC48667441ABE357563C8C6A610672B509377D9AC",
		INIT_04 => x"D08AE2719BE3EB78AA7CE3D2A5D72F4E77D01C44006B03B6C4133519524D1988",
		INIT_05 => x"B7D5D9BCFB1495690F86EF4DF2985B68EE56E631DF8B27B0F8833715C29155B9",
		INIT_06 => x"488DD52630FF1269E8361554750BF7DFC048B4975C114767C927F5AA63AD6AF4",
		INIT_07 => x"4F68B227F953E5CC6E55864E573F0FB4D8FC496206E8CADE2396FEDA4DB6D8A1",
		INIT_08 => x"0888A53B152261D32623CA060D9EDED1BD2100CCA2F899F56517E3D946C07991",
		INIT_09 => x"D1323D298760A0C630E1A02B84C7DCF2D0B14C918E098D0937830E356BDE216F",
		INIT_0A => x"487F81EC153B255CC00E9D8385371328B3D45349A3DC698BB86736F802FCD921",
		INIT_0B => x"3D76A4DEFC3E0FA3F9F4DEDF7C553C6FE61CD85EECBD621408223252D8EEE9C5",
		INIT_0C => x"4D86EA8503E72E4897A31E1A4235EABAC9ED5959F2AC3513B2AEFF6655B84F0C",
		INIT_0D => x"E39E8623ECED06B79A887BB666F86CCB2D1407968260AF6B35AC1644C7F1799D",
		INIT_0E => x"A51744CA0292B20E21D5E546E436C1619F3EDC4B1E82F6A78548A773F12FBB1D",
		INIT_0F => x"983D58E4184DAF4D83C69B445D573BB6333F967769BF5FBD7A2149E8AFF1DEDD",
		INIT_10 => x"16EA4DE6C8400495385CBD57A0DDC0CB41C3BA558289339633C15CA70FEA1FB4",
		INIT_11 => x"F9B2CD5AD0D67259DC33C1763AA02C4F1C44617D86B1DB9035E2D2B7B98A4DD4",
		INIT_12 => x"812380E1A2719C990E54E220E1F064EC49F703FEBDB4E24E02806D41BC0B0AC8",
		INIT_13 => x"4EC4C02431B130D3CA06E72E446216DEDB3C160C9EA93C853B2250A8C435852B",
		INIT_14 => x"CC2B3FFB4C4B1FA89EDD288F5DE85F99451883524231CA19AD3656CD247DA427",
		INIT_15 => x"00B9A76378E819C2F813ACBF2BD5469ACE0424DA6991A60F66CF3FB93551ABCC",
		INIT_16 => x"6E23FB123D87AD848EBBD1729792B743DFC94FA3DF4AFE3B5FA9804D17CDE843",
		INIT_17 => x"0540148B6827EA3E82F255C60108D04B6CE5BE9A53115AD26563C3E7C97B1294",
		INIT_18 => x"6E43D63C222AE3BE2E8EED6D90CDC0920697DB13F55892EFAF88FBE5E6AF2891",
		INIT_19 => x"3BFB1DFB64EA8588693EB4B85B963B5E92762E963F1633940FFCF858281C4A82",
		INIT_1A => x"189C9010A53535A4423B5C15C47D0C1DCE20A6EC4727C4E32ECA126B81872E55",
		INIT_1B => x"B53FED5185A8709C4B0CBB0F4C75AA9BADE0BE715340D7E79E8A300C40BF4FD3",
		INIT_1C => x"0446ADE103691EECEDAA5C33E64DB252942B7F756539C7EE8C68D7E593829A87",
		INIT_1D => x"541D0105007819A37B94ACD451AD0627D45C66E45F137E5FB8CF4B5BDD124690",
		INIT_1E => x"CA2F6FB5DC7A6D5A7B5315A374C24A3544713B0741DA3E336CA646D34D69D2EE",
		INIT_1F => x"A4EA0B304DF5BC15287C2A7DDB1CDB4F199004F415AAA5FF757BDDA714A4030B",
		INIT_20 => x"1F80BB4B2699CA6C0EE3C94303FD075F5D8E624413BF65380732F7794BD70C1A",
		INIT_21 => x"C793ABBCAA05250F0F93C5241198585F10A8DE6B07F58E1FB524E6808704F597",
		INIT_22 => x"50E763251C317C7AEBC978AE68627AFB3209FA5F02144D8067FA912271A5409F",
		INIT_23 => x"EB6680DCAA04568290D5441C016723CD2C6D8D45158D6B0C5C31B2D587522EA3",
		INIT_24 => x"8B02096A46AF96B6D77B745A4F25BE8C0883BBA81736C25C597739FCA219EAA8",
		INIT_25 => x"D5275D415F3E07E2EFD03A5181BD3D30F7CA40BA212E280623B56A632037F62B",
		INIT_26 => x"FA4FEDBFB98B28E5B26747489503D7A240C7EA5D65435E0F581544D73D6E4155",
		INIT_27 => x"05057B0F8E7A56E03D9C1D39115ACF8F122AA8753FBCCD69BBC9DA89DCEA6288",
		INIT_28 => x"9E9D4F2E6A0FA074089A76258BDAC59565D8C4559CECD61AB351A24FD652AB8A",
		INIT_29 => x"98B7B8625573C386AC28D5099F17B432FBA03A3DF5F0D4FECB878325D8D040F5",
		INIT_2A => x"C2842FEC2C5C8CFF8247937ED20B4875D88BCE5A094C50BD5415C340B9973BAC",
		INIT_2B => x"5174F4DE971ED9175653CDC84E45E5978CA4DB481E4D3E7F406CA3C7E062D3A6",
		INIT_2C => x"DAAAC5CEA75D57A81E442D53E2EA8DDA30C38608502E232E8B07773E39964F55",
		INIT_2D => x"57AAA5C361C909BC0E8D20D7C7249B03178706DD527F69183B1205E98FF987B3",
		INIT_2E => x"64715F6A3E8D268CB92061AC2398489B6F2348367D18C26E5780D24690DAEA45",
		INIT_2F => x"44587CDDC45C91E1A2CA7AEDC95603D31C446C728956770986F57D4927D15C32",
		INIT_30 => x"EC5065063A42A1184004D9B78C102353E5653715B52722167B670C345A9E286C",
		INIT_31 => x"4D2436A7985F3EC4F564D7A2C5DF03D75DB62703812B9CBF42717D0FCD528C3C",
		INIT_32 => x"00DE1C278B0EF98237595B9D27E4EE67177DE6653FA2885A3B74CA66CF45478A",
		INIT_33 => x"C52B981DB25CF31AD9D6E72D3BFFC736EE507E065D0FF53778738636CD353B30",
		INIT_34 => x"4E59124EB038A30327BD74252FBA8CB4775774C2FA2DA73647B5B59FAB63AF43",
		INIT_35 => x"E1048E141235BB66B172AC58FB722F02F8B151EBF64A04578AECF347C29A400D",
		INIT_36 => x"E1950BEC0E0A344DF58A461826FD237E0CBA08364C4825780B3DC832DD184B68",
		INIT_37 => x"D3BD115A719569FC8CADDE3BB759D98114690B8D6A94FF3CE7E703D9448C0CDF",
		INIT_38 => x"BB117345FE411E664279B3269F78BC9D6630A1F731057E82086175744831E72C",
		INIT_39 => x"6DABF8058BD20E4EAD1BED828D422D4AB0A10AA5C39C2C3A07FD945C1BAC4837",
		INIT_3A => x"708DD6B86A4767889AA6D54922D525A9B2952D71C85982253232FC6B2DD68E56",
		INIT_3B => x"D92608B2E8AB73ECBD1B6ECB280DE2F4629D649B006F6BD473071734BA1DAED3",
		INIT_3C => x"91F8CCCD7EBEBF8E6EFEB808B4AC38DBDAC8333A178AED3B17EF9DD6504B3F89",
		INIT_3D => x"286D5D152E50D42086473C0B51DAFE0C7BD6D3CAE4BC7611C4955C80F0029B18",
		INIT_3E => x"CBE66E2BF17781BE0E76458EF24A0C97CDDA7DAA7CA3E9D9AD9902B3DC41C65A",
		INIT_3F => x"11111111111111111111111111111111BCBC97CFC194CDCC6809281D370204FF"
	)port map (
		DO   => doutout,			-- Port 16-bit Data Output
		DOP  => open,				-- Port 2-bit Parity Output
		ADDR => addrin,				-- Port 10-bit Address Input
		CLK  => clkin, 				-- Port Clock
		DI   => (others => '0'),	-- Port 16-bit Data Input
		DIP  => (others => '0'),	-- Port 2-bit parity Input
		EN   => '1',				-- Port RAM Enable Input
		SSR  => '0',				-- Port Synchronous Set/Reset Input
		WE   => '0'					-- Port Write Enable Input
	);
	-- End of FRAME0002_RAMB07 instantiation

end FRAME0002_B3;