--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
--	Grupo de Apoio ao Projeto de Hardware  - GAPH
--	Projeto X10GiGA - FINEP/PUCRS/TERACOM
--
--	M�dulo:	Mem�ria - Gerador de Frames - Prototipa��o
--	Autor:	Jeferson Camargo de Oliveira
--
-- 	FRAME:	0003
-- 	RAMB:	00
-- 	CONJ:	B
--
--	M�dulo gerado em 17 de July de 2008 �s 16h55min pelo
--	programa gerador de frames OTN do projeto X10GiGA.
--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

----Pragma translate_off
library unisim ;
use unisim.vcomponents.all ;
----Pragma translate_on

entity FRAME0003_B0 is
port(
		addr	: in  std_logic_vector(9 downto 0);	-- Barramento de endere�os da porta
		clk		: in  std_logic;					-- Entrada de clock para a porta
		dout	: out std_logic_vector(15 downto 0)	-- Sa�da de dados da porta
	);
end FRAME0003_B0;

architecture FRAME0003_B0 of FRAME0003_B0 is

	signal addrin	: std_logic_vector(9 downto 0);
	signal clkin	: std_logic;
	signal doutout	: std_logic_vector(15 downto 0);

	component RAMB16_S18 is
	generic(
		WRITE_MODE : string;
		INIT_00,INIT_01,INIT_02,INIT_03,INIT_04,INIT_05,INIT_06,INIT_07,
		INIT_08,INIT_09,INIT_0A,INIT_0B,INIT_0C,INIT_0D,INIT_0E,INIT_0F,
		INIT_10,INIT_11,INIT_12,INIT_13,INIT_14,INIT_15,INIT_16,INIT_17,
		INIT_18,INIT_19,INIT_1A,INIT_1B,INIT_1C,INIT_1D,INIT_1E,INIT_1F,
		INIT_20,INIT_21,INIT_22,INIT_23,INIT_24,INIT_25,INIT_26,INIT_27,
		INIT_28,INIT_29,INIT_2A,INIT_2B,INIT_2C,INIT_2D,INIT_2E,INIT_2F,
		INIT_30,INIT_31,INIT_32,INIT_33,INIT_34,INIT_35,INIT_36,INIT_37,
		INIT_38,INIT_39,INIT_3A,INIT_3B,INIT_3C,INIT_3D,INIT_3E,INIT_3F : bit_vector
	);
	port(
		DO   : out std_logic_vector(15 downto 0);	-- Port 16-bit Data Output
		DOP  : out std_logic_vector(1  downto 0);	-- Port 2-bit Parity Output
		ADDR : in  std_logic_vector(9  downto 0); 	-- Port 10-bit Address Input
		CLK  : in  std_logic;			 			-- Port Clock
		DI   : in  std_logic_vector(15 downto 0); 	-- Port 16-bit Data Input
		DIP  : in  std_logic_vector(1  downto 0); 	-- Port 2-bit parity Input
		EN   : in  std_logic;			 			-- Port RAM Enable Input
		SSR  : in  std_logic;			 			-- Port Synchronous Set/Reset Input
		WE   : in  std_logic			 			-- Port Write Enable Input
	);
	end component;

begin

	addrin <= addr;
	clkin  <= clk;
	dout   <= doutout;

	-- FRAME0003_RAMB04 instantiation
	FRAME0003_RAMB04 : RAMB16_S18
	generic map (

		-- The following generics are only necessary if you wish to change the default behavior.
		WRITE_MODE => "NO_CHANGE", 	-- WRITE_FIRST, READ_FIRST or NO_CHANGE

		-- The following generic INIT_xx declarations are only necessary
		-- if you wish to change the initial contents of the RAM to anything
		-- other than all zero's.
		INIT_00 => x"C23CFF00EF967228CE2CF081732D544674AEAE47E4DC39073435925DF3FF1706",
		INIT_01 => x"53282FE2E4D839C5E873A210EFF194748B4CA6FF63FA5FE54CCB7E88E4B49C69",
		INIT_02 => x"ED0BE7AD8745D71C52A340DD07D8C144028C2E4ED45B4DF8CE76ED3F1E0C5391",
		INIT_03 => x"D3FE87469B63858FEE3EF576F6027A8933B89CCACBB0E5FBA940D2AB7DB4C7FD",
		INIT_04 => x"61E47D35BCE779E0A6F8823F2C7B1C13E854E38BE484B0E85E88A25121FDF41E",
		INIT_05 => x"255717A609519A8D066862B48535FD90080766B1C57A273C82A4985670A16A0A",
		INIT_06 => x"E9406ED17DF6BAFE461C1B2541FB39BFC46C8B1E8DFE0164AC1661984080CA74",
		INIT_07 => x"FE05453442F18DAD32CDBBB4D5F1567E297A2FB5B14FE3A30366C77364AA8ECE",
		INIT_08 => x"254C10A4AF5C5C8B84645F92A8E03A84A5AEA9D85D7D170E6AD68C7BAE1AE0FB",
		INIT_09 => x"B8254D45F321D7F26FD7B1685A3AB6639FDD5977568A6E1143E7F1606E73A65B",
		INIT_0A => x"5A50CB8EB44BC1E01B3940617CC60A05E1930BF289EF9672EF8CC6923315E67B",
		INIT_0B => x"5B4114D29E4B0848C6DF7125FA58A930D3B8B85D749E80527898ECE48723BAC9",
		INIT_0C => x"60E3735CE2FBCED2BD56C535977E2F5AF915FAF70C73EC304AE452836A04DD1C",
		INIT_0D => x"C873476EB9D134E6DCFF8FAB9E865D7A05504116A0F4E1FCEF518B2293327B08",
		INIT_0E => x"62FBB86564F313BA8947E71642E56967DE60BE16E49592B552C40A05FFFA123B",
		INIT_0F => x"5313D4C001145EEB9B93A50E19AE232E2B865B078D8197A13CC40869A87CCCEB",
		INIT_10 => x"7DFA3DFC98DD4AA799856ECF83E0B0B1D79DD1BAB6A77FE8B97A3589040A3BFE",
		INIT_11 => x"7745DF428C35DC079EFEF1C1D4C2D294037D9D5FEDC1DCA73C12BFD654A1E918",
		INIT_12 => x"59941457C87278E867DC5BBEEB913532FFB89287C28824166526AE37FC1662EF",
		INIT_13 => x"68DFF17F27C42294DD204995E906DB6ADA5A11762CECF05A07E644678A4ABDAE",
		INIT_14 => x"44FEEF861AFCEBA8E108CA7437ACE158FAED71250FB64B5D76C6E206ECC9F576",
		INIT_15 => x"7858834250E361C1B6D23745A182FBB0FB383B8D6D57BE082C603FFED91D6B2A",
		INIT_16 => x"BC9B7A99605C772831AFF76D08D39730E24E70A3A1CB6843C713F541EB818C59",
		INIT_17 => x"6D1643248E85AF6D0B82E5F9625756AF1ED0DCBDF8ADD995F23674C0B278D46F",
		INIT_18 => x"28298C5FD230AFD24CB2FED2287EDBB4E3FB0755AAFD5966C54DF044C9682730",
		INIT_19 => x"C869EC141F229D2288F1A0BD30B769CA41903E3969CB909E9AF7C68E3F20B6AD",
		INIT_1A => x"7EA3C97C4E5E6A757FDD3E1F28A560ECA1149066AC32F0CC51B0893F3A5D27A0",
		INIT_1B => x"8D97B0528E61BD8539C774CA356532819EED281A8FD8AFFE3763FF325DBE0A60",
		INIT_1C => x"706F3D73EBE219318D7DD8EB337CB88DD376EF04393F1893A3AE1475DD8E4EB5",
		INIT_1D => x"339A4F3B3F025C75E5A9A6A2C576BDDEEF32E699ED5C0448A785613A1C9D66D9",
		INIT_1E => x"2CC19A024E122792FC832BD96C60689371A568A8D14F15C6574FF4FAE8D3AC50",
		INIT_1F => x"A1B4AE24BACD3557DB7446E126BB6C24FEFDE1187D8AD3249C54AAACBD0F62EC",
		INIT_20 => x"C6BDA16083311F5FCACA4E2916FB434DE1DAAA8DE02C8E1125ACA2102C82CB24",
		INIT_21 => x"F3B68E3E7CF6191EBB35202EE3DE24AA11E122CC39F8B18A5564953F4A89C154",
		INIT_22 => x"B4D20991EC68266E433903D90898B088CC5CA4BF0FF55405386C9A609C771FED",
		INIT_23 => x"C1594D4839D33324588BE3D7AEDA1452A84CE9A1D8853B9FF489CC28ABCB9530",
		INIT_24 => x"95F40DC5443E643FD73012C7A1B1E8DCFB41A6C1AC5A30E8B0825840654BD2F9",
		INIT_25 => x"F8F18A7CF044C99392910965CCC8FC8521E8A8C8D35C8579455CA77765716BF6",
		INIT_26 => x"753BA276A108AF11657F504F24F9176D3DDAFA3E5267FDDAB3A18BC950C75540",
		INIT_27 => x"5E5887F4B0D2B817F3180F364CE50A947A7FAD0A2C15DFDA99304354C8E7E048",
		INIT_28 => x"F7C0F83D1B3144F7974BC1C7A3C0D63548FAABA5156D340A66AEF74363028915",
		INIT_29 => x"8602404FC7E91B2B696E49B150941DCA15041B76CECC1BC4D86DB06C5D41D920",
		INIT_2A => x"5577C6866796A1F6CE9743B3638E8CC3944EBD2BAAC537D40BEB3814A46D63E1",
		INIT_2B => x"08FBD4E96D1123AC1535D019D002F65B533DA292B92176430E902B3ADEED954E",
		INIT_2C => x"48BFAF10394E345BFDEAF3C9B70EE25424D7F2AE55331BCE540293132B6D93D3",
		INIT_2D => x"FE61E94AEA64EEE94373DC368A57F06E3E39263D39DDE09EF3F26644869F3502",
		INIT_2E => x"F43AB1972F6C01D3E315F205E3F250AA33128177A2A73DE1EEE3BC78BCAC4641",
		INIT_2F => x"187C81C03DD07048B46CE75028F716129494C8BA907ECB2DB6EFD71C87F5A501",
		INIT_30 => x"AB20DC382F5EF274607C527FF3ABBC7F8D699533386D883581E2491413290842",
		INIT_31 => x"44A083B7C72B14EDE572B809295E2F001B1109F6C8DE79A514C1196CA909BD29",
		INIT_32 => x"3ABA773F2B43311DA05532B428EA14012E1D9BD32A0D4655B718DA58385C905B",
		INIT_33 => x"B5C5936B3A0DAAD73C5FA5D8E22491DD307ADD9249266926EF71799C8E76678E",
		INIT_34 => x"3E803D2181C237BA06BB76BED26532EB4C133E0EF70F65A7F6E7F0E09894E0D0",
		INIT_35 => x"F45C67D6C58F9A06249EE2D7703A56271A711BE037CEBDBDCCBBD87B684022DB",
		INIT_36 => x"6E8D8158C1C8C754E3E35A17457CCFD2F9A5218564DDE4797B0866051B566257",
		INIT_37 => x"99DAAE36AC1C03E2EEBB08B9C46C7D8781078B527D8B05A426988531085CA465",
		INIT_38 => x"E42364F7759C2DC1A2A7C0C2554EE907575DC1B2AA1DE71EB309596EA31683F1",
		INIT_39 => x"0D3596A4269588491F26E7710B7FE2B0DF20A4D5E902B861372B7CCE7AE2CCBD",
		INIT_3A => x"6CABE7A330ACD418F016950E848E2B2E331DE438D5ECE91BF591E968EEFBAA5C",
		INIT_3B => x"CF7AE7C7612A9927A0F9542DE5CA47899797CE491E06D1D59B82758B6B2A9674",
		INIT_3C => x"03F1F755D33BCEBFA60842BA28C0F3701F83CC1406CDCAF8E4B996113CF71A96",
		INIT_3D => x"E49629AC99D950EA0DEDA2502F918AD600AAC1F04CDE2C41453E126C0F4F9D3B",
		INIT_3E => x"05F5A1967AA0B1CC34F8CF04FEE27D5CAABF8EAB68F01970060ABFB1682138C6",
		INIT_3F => x"11111111111111111111111111111111DF12CE54982EA3903417081D73551319"
	)port map (
		DO   => doutout,			-- Port 16-bit Data Output
		DOP  => open,				-- Port 2-bit Parity Output
		ADDR => addrin,				-- Port 10-bit Address Input
		CLK  => clkin, 				-- Port Clock
		DI   => (others => '0'),	-- Port 16-bit Data Input
		DIP  => (others => '0'),	-- Port 2-bit parity Input
		EN   => '1',				-- Port RAM Enable Input
		SSR  => '0',				-- Port Synchronous Set/Reset Input
		WE   => '0'					-- Port Write Enable Input
	);
	-- End of FRAME0003_RAMB04 instantiation

end FRAME0003_B0;