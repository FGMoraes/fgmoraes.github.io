--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
--	Grupo de Apoio ao Projeto de Hardware  - GAPH
--	Projeto X10GiGA - FINEP/PUCRS/TERACOM
--
--	M�dulo:	Mem�ria - Gerador de Frames - Prototipa��o
--	Autor:	Jeferson Camargo de Oliveira
--
-- 	FRAME:	0001
-- 	RAMB:	02
-- 	CONJ:	A
--
--	M�dulo gerado em 17 de July de 2008 �s 16h55min pelo
--	programa gerador de frames OTN do projeto X10GiGA.
--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

----Pragma translate_off
library unisim ;
use unisim.vcomponents.all ;
----Pragma translate_on

entity FRAME0001_A2 is
port(
		addr	: in  std_logic_vector(9 downto 0);	-- Barramento de endere�os da porta
		clk		: in  std_logic;					-- Entrada de clock para a porta
		dout	: out std_logic_vector(15 downto 0)	-- Sa�da de dados da porta
	);
end FRAME0001_A2;

architecture FRAME0001_A2 of FRAME0001_A2 is

	signal addrin	: std_logic_vector(9 downto 0);
	signal clkin	: std_logic;
	signal doutout	: std_logic_vector(15 downto 0);

	component RAMB16_S18 is
	generic(
		WRITE_MODE : string;
		INIT_00,INIT_01,INIT_02,INIT_03,INIT_04,INIT_05,INIT_06,INIT_07,
		INIT_08,INIT_09,INIT_0A,INIT_0B,INIT_0C,INIT_0D,INIT_0E,INIT_0F,
		INIT_10,INIT_11,INIT_12,INIT_13,INIT_14,INIT_15,INIT_16,INIT_17,
		INIT_18,INIT_19,INIT_1A,INIT_1B,INIT_1C,INIT_1D,INIT_1E,INIT_1F,
		INIT_20,INIT_21,INIT_22,INIT_23,INIT_24,INIT_25,INIT_26,INIT_27,
		INIT_28,INIT_29,INIT_2A,INIT_2B,INIT_2C,INIT_2D,INIT_2E,INIT_2F,
		INIT_30,INIT_31,INIT_32,INIT_33,INIT_34,INIT_35,INIT_36,INIT_37,
		INIT_38,INIT_39,INIT_3A,INIT_3B,INIT_3C,INIT_3D,INIT_3E,INIT_3F : bit_vector
	);
	port(
		DO   : out std_logic_vector(15 downto 0);	-- Port 16-bit Data Output
		DOP  : out std_logic_vector(1  downto 0);	-- Port 2-bit Parity Output
		ADDR : in  std_logic_vector(9  downto 0); 	-- Port 10-bit Address Input
		CLK  : in  std_logic;			 			-- Port Clock
		DI   : in  std_logic_vector(15 downto 0); 	-- Port 16-bit Data Input
		DIP  : in  std_logic_vector(1  downto 0); 	-- Port 2-bit parity Input
		EN   : in  std_logic;			 			-- Port RAM Enable Input
		SSR  : in  std_logic;			 			-- Port Synchronous Set/Reset Input
		WE   : in  std_logic			 			-- Port Write Enable Input
	);
	end component;

begin

	addrin <= addr;
	clkin  <= clk;
	dout   <= doutout;

	-- FRAME0001_RAMB02 instantiation
	FRAME0001_RAMB02 : RAMB16_S18
	generic map (

		-- The following generics are only necessary if you wish to change the default behavior.
		WRITE_MODE => "NO_CHANGE", 	-- WRITE_FIRST, READ_FIRST or NO_CHANGE

		-- The following generic INIT_xx declarations are only necessary
		-- if you wish to change the initial contents of the RAM to anything
		-- other than all zero's.
		INIT_00 => x"5B29EC447D921EEC6C1BE0E241B83B9CF11BC1B717C49551E8D187C1131F2828",
		INIT_01 => x"FE1FF449BD40E58BDF4907CDB9BA24D77252F22077BC542489BFCF1DBE34BD7A",
		INIT_02 => x"5680BF9F37845B534A5DC541BCB724035AD3148D82F50AED0087F5A9B0BF577D",
		INIT_03 => x"771C81B981AEF4C656E4BD059FDCDE37C81B81EACB5CB9530B45425B4F55934D",
		INIT_04 => x"4C63B99DFAD61C52606E02EE208A80C24AA08619C3BC4F18AEDFF2C07060E06D",
		INIT_05 => x"807BC205EED94C66E6A96F97933945B6785F681CEA074AF33A240A80B7C0D135",
		INIT_06 => x"E682F5109D20BD9C30E54FF694B3C0AE63411F167F04CCB36C2C23DC1896F804",
		INIT_07 => x"CE0A1B0D73E930BF362D11275001EAA2CC5788A888CF8B8ED1811699A4698F5C",
		INIT_08 => x"96EAE9937E67302F1FA12EE2A963DC744F63E70B63176DFFD5C756CD05F05538",
		INIT_09 => x"E29BEB5AE30A6CE9DCCF6466C2CB71B16A296ADDB027946F6268F21596B10524",
		INIT_0A => x"70494A851623B2B8EEDB0A663A78DC5C45D544E67F951D59B46D43A058C17B60",
		INIT_0B => x"A5EC35B15E92D269EDA74FD1C4DBF2E266D2215F5ED45184A57672011E98D92B",
		INIT_0C => x"4260D8DD714E4029F253CDEC04C9DCBABB9F30BDB286FF0928DC871B99B4A811",
		INIT_0D => x"25923A630184D57F2A81B72738F6F3403167BA5DA31B095B7BFDD972D0804DB2",
		INIT_0E => x"1DF75C2A384550FA5DFF30D244A229D579132EE807F861A9BAE79E8796D464CD",
		INIT_0F => x"BBB77D37CFFD70E201B2D2B96134D430269E90A448F00281C17A3756D225370B",
		INIT_10 => x"0247E908E693CFFD280B66BC0D18BA7E9BD650F0C1D5FFDEF8955D65FF142DF2",
		INIT_11 => x"870EE836F13B44D904E183277B73B71E97A0426890F2E8D221C0CFD213CA4942",
		INIT_12 => x"F3F5DD683B4CD7D96865652BBFB9AEEB0A8E00AF69DD5C51458FFE9A2567FAC8",
		INIT_13 => x"0756A4A5A4E4B0EFEB39840EFDABF294EC8EF4B089152EDA5F9781DB6DF6CB97",
		INIT_14 => x"DD412721638593F8F42FBCC32F52623D6AE0EF26A723CB52B19C74A1B004EA60",
		INIT_15 => x"B1C3506DA21B5485D7650164A1538455CF3F6E4786A26FFE5806DCF975C39458",
		INIT_16 => x"FEF7EE67415ABF8949837394BC07390B02C16877D09EF9802B9EB06D936615FC",
		INIT_17 => x"16B0CE8F00328836B2B9B2E7E0190636AB0975D4460CD1D784D57D6E6BAA71F9",
		INIT_18 => x"03793AA9C51CE4FDB67547EF562977EA70BA85B3820F5F7FD373900F236AA402",
		INIT_19 => x"3BCB4DA9430480CD170C0C662BAC5C6AF03F423CC3B8C303D744B10459166261",
		INIT_1A => x"384A8A94C5180110B679EAC46ADEBEB7FE53EB148C795751F6CBEA9F6AD47061",
		INIT_1B => x"DF9CFD948ECEFC17A53758CC5A83F70A56977AA6694A473254F7597C4732C160",
		INIT_1C => x"C67DF8FE4E01862A7E85A4ABFBA143D9D3EE235593A1266E0498F5002E26A029",
		INIT_1D => x"9A7D5147A5EEB86D1EE781BAA986FC149A29B66908BF7C7A30B979DB1D8A63AD",
		INIT_1E => x"67AD589F582E8676431BB00F8E61AB8AFCCEF9A56D3D4819FA2FAEADE9666505",
		INIT_1F => x"DCB1CB43B6B497F16189101D92A1200FB81E8BEF6956835C4B54E78D02BDC815",
		INIT_20 => x"9972AD93F9C83F47AC0E920287E62E90D3C0FF9CC35F6DD0277D10893602A5BC",
		INIT_21 => x"494A236FFF4744811FD859653D83629BDF10FB1238C75983BA6177594FCDCFEA",
		INIT_22 => x"E9C2C7BEF923F7F8145ECF2320CFD9C9DB69C3079A2532AD098A7D57C1B4A019",
		INIT_23 => x"68CCB0DC4EDF1067CB428F0085D754709CDE87795F24FA21EDC40DF3FCA392AA",
		INIT_24 => x"A8DE28121AFDFECF3C9954629BEA240BDB5E89166970DB6638DC10EF6154F8C7",
		INIT_25 => x"966E607059563EE509CE568BAC72A4C53C343894FA0298D97AC213A174564CDC",
		INIT_26 => x"B7321CB6B0CCFB4D5D975C3DA0D297FBB7A4013FB63070CE7151943A9F4073E9",
		INIT_27 => x"C1801BF014DB6802E262D86A3FF25367BAD39027888872046BE225031AC31692",
		INIT_28 => x"070014DD57D5CEA8DBA184A9D4F9014E445A5D621E366721AD927672076A25E6",
		INIT_29 => x"134A2D465DEBBBA5FEDA08907B4BC5E5F824AB8335ECAF7080234E8122849C57",
		INIT_2A => x"FB9C2CBCF9EB496D9C2DDF365E30B8D82909A0D749462AE7DAD2210E78E99F1F",
		INIT_2B => x"396CD93DB6E1D9B20485DEF8679B1E6CC55165371A6147500ADC0CAB371B687D",
		INIT_2C => x"72219F9F4C6C877A516727D996708540FB340CB73D96A17C51A1698F34847A84",
		INIT_2D => x"261FDAB1CFE7130AA088FE8E454EA077994F9E85486FB5AA0BEDEB36EF457B70",
		INIT_2E => x"C549527949DC73F5C35B78E990992B80CAD378167AF676F8ADAD7A6B7CA24357",
		INIT_2F => x"25257FFCF30D7D67E39D1FD366ECA95B2DD61CB8F68690355C191AE19F797F29",
		INIT_30 => x"7D7299840F06B194EE85A91D3F7A6107C6CD0CDD61B459CBD6301B4385C560B5",
		INIT_31 => x"EE676DA53EFB5460CF004D029B5D746E9A7E51094DA179A8C59D61136EC03104",
		INIT_32 => x"C2E24AEB4FDF16D01C4F130299C80C0AEDF22EFC607ABED989BC3505563DD63E",
		INIT_33 => x"17D148F3C11F43B5A4C558C6BD479909BEF5509CF2F6E4DEFB933D4658C353D7",
		INIT_34 => x"1D7C3B40A0058D1C6A5E2FC97D938F5C50EF2E646B6FAA418C7C815BDCC801E5",
		INIT_35 => x"11648D4284C0D53549168A27BE7036395B42AB84DEE27F8E58DD93525A3924D3",
		INIT_36 => x"32A9D704FEA9FFAC621C15670CCF924AE5CCC32D53FCBCA7BAAE0653CCBE8966",
		INIT_37 => x"D25498DE75FC10B46729FC75AB40AAB22EEFDAF8B869231A50578630A7DB7A9C",
		INIT_38 => x"7A4BE55E6066AB4B0B3A0AD0177146A35010D60B5528FD939EC151F4AB964E07",
		INIT_39 => x"BCE9AE4D8B5353645289CB4A79150B03C76CFDAFE7BAB9C3E6656C3C24BBA3B5",
		INIT_3A => x"CF1F237D69388CE4627E333BFA0ACE081587D17D5DB0D55BB503611791A971AB",
		INIT_3B => x"A57101C40274AC78BD8D7F7CCA66CF3FCBCC36FCA3F87721F56CBDB5C1BD7996",
		INIT_3C => x"606A3E58FACC60824041FA51C93E1400A488C3D591B3AB5C378F5D5AE577CBA8",
		INIT_3D => x"9B87632832C971FAE6B2AFB1B73A84DFB292E93A36DBC28EDD84A914C5750192",
		INIT_3E => x"DD58B75DB470DC5056A0FEF7A17DAD56904FA22D2B722FBDDBC1DAE41B52E978",
		INIT_3F => x"08A2EBC79BE9CF0FC2D5C49FF4AF2674395F44731AD0132E6045EB5B0F83BB3A"
	)port map (
		DO   => doutout,			-- Port 16-bit Data Output
		DOP  => open,				-- Port 2-bit Parity Output
		ADDR => addrin,				-- Port 10-bit Address Input
		CLK  => clkin, 				-- Port Clock
		DI   => (others => '0'),	-- Port 16-bit Data Input
		DIP  => (others => '0'),	-- Port 2-bit parity Input
		EN   => '1',				-- Port RAM Enable Input
		SSR  => '0',				-- Port Synchronous Set/Reset Input
		WE   => '0'					-- Port Write Enable Input
	);
	-- End of FRAME0001_RAMB02 instantiation

end FRAME0001_A2;