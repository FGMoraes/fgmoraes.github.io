--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
--	Grupo de Apoio ao Projeto de Hardware  - GAPH
--	Projeto X10GiGA - FINEP/PUCRS/TERACOM
--
--	M�dulo:	Mem�ria - Gerador de Frames - Prototipa��o
--	Autor:	Jeferson Camargo de Oliveira
--
-- 	FRAME:	0000
-- 	RAMB:	01
-- 	CONJ:	A
--
--	M�dulo gerado em 17 de July de 2008 �s 16h55min pelo
--	programa gerador de frames OTN do projeto X10GiGA.
--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

----Pragma translate_off
library unisim ;
use unisim.vcomponents.all ;
----Pragma translate_on

entity FRAME0000_A1 is
port(
		addr	: in  std_logic_vector(9 downto 0);	-- Barramento de endere�os da porta
		clk		: in  std_logic;					-- Entrada de clock para a porta
		dout	: out std_logic_vector(15 downto 0)	-- Sa�da de dados da porta
	);
end FRAME0000_A1;

architecture FRAME0000_A1 of FRAME0000_A1 is

	signal addrin	: std_logic_vector(9 downto 0);
	signal clkin	: std_logic;
	signal doutout	: std_logic_vector(15 downto 0);

	component RAMB16_S18 is
	generic(
		WRITE_MODE : string;
		INIT_00,INIT_01,INIT_02,INIT_03,INIT_04,INIT_05,INIT_06,INIT_07,
		INIT_08,INIT_09,INIT_0A,INIT_0B,INIT_0C,INIT_0D,INIT_0E,INIT_0F,
		INIT_10,INIT_11,INIT_12,INIT_13,INIT_14,INIT_15,INIT_16,INIT_17,
		INIT_18,INIT_19,INIT_1A,INIT_1B,INIT_1C,INIT_1D,INIT_1E,INIT_1F,
		INIT_20,INIT_21,INIT_22,INIT_23,INIT_24,INIT_25,INIT_26,INIT_27,
		INIT_28,INIT_29,INIT_2A,INIT_2B,INIT_2C,INIT_2D,INIT_2E,INIT_2F,
		INIT_30,INIT_31,INIT_32,INIT_33,INIT_34,INIT_35,INIT_36,INIT_37,
		INIT_38,INIT_39,INIT_3A,INIT_3B,INIT_3C,INIT_3D,INIT_3E,INIT_3F : bit_vector
	);
	port(
		DO   : out std_logic_vector(15 downto 0);	-- Port 16-bit Data Output
		DOP  : out std_logic_vector(1  downto 0);	-- Port 2-bit Parity Output
		ADDR : in  std_logic_vector(9  downto 0); 	-- Port 10-bit Address Input
		CLK  : in  std_logic;			 			-- Port Clock
		DI   : in  std_logic_vector(15 downto 0); 	-- Port 16-bit Data Input
		DIP  : in  std_logic_vector(1  downto 0); 	-- Port 2-bit parity Input
		EN   : in  std_logic;			 			-- Port RAM Enable Input
		SSR  : in  std_logic;			 			-- Port Synchronous Set/Reset Input
		WE   : in  std_logic			 			-- Port Write Enable Input
	);
	end component;

begin

	addrin <= addr;
	clkin  <= clk;
	dout   <= doutout;

	-- FRAME0000_RAMB01 instantiation
	FRAME0000_RAMB01 : RAMB16_S18
	generic map (

		-- The following generics are only necessary if you wish to change the default behavior.
		WRITE_MODE => "NO_CHANGE", 	-- WRITE_FIRST, READ_FIRST or NO_CHANGE

		-- The following generic INIT_xx declarations are only necessary
		-- if you wish to change the initial contents of the RAM to anything
		-- other than all zero's.
		INIT_00 => x"59B4866944E3B37B74317646431C4D6F0F0C7AA5D5F77DCABD54D2CE05D2F628",
		INIT_01 => x"2C533DB8162DD2E0C06ED476F0123DC0C179FE337E8383436BBDA63E9AF0FAA2",
		INIT_02 => x"F9375939F4E5ABE74EBBBD482896E1FD4BC78FEDE79B6DA1B4D5792E4285B331",
		INIT_03 => x"FD17CE3819283BB68E624667F85B58164FF1E452AECFBBF349918B57CE69AAB8",
		INIT_04 => x"1C870445E390D224C10296C0EA2E6E9758FA83736E6C68DFDE2FE817B2847F76",
		INIT_05 => x"3C1EB38EBA6D2F7498DB9B82C074F573685D34CCF604CE77C9079E7F446E9F0A",
		INIT_06 => x"6A09D72D3B94F5E8A03F4C19548BDBD1CF9E79AF5138D1B817177526994EED14",
		INIT_07 => x"2B75E646DA00C5EF3FA2216D0BAC81FD26EDCAB94EAD0312FE024C948A27FAF6",
		INIT_08 => x"877E49FEC2697021EE8E89FDC4A4B72D8FDEB563A48286DDBD18E4964CB99FE1",
		INIT_09 => x"DF1515A08CDE89F3855E0B7667FF6DCB1C4FA6AC60D1C495D52D2EE7A7975E28",
		INIT_0A => x"F4DB3C04E2B0E3E0ACA7A4C55FC571AC960EDB48979C9516133CB5B4696C563D",
		INIT_0B => x"5194E63CD60453E0FD174A68E5CC418C8B498723EC83114E6D7E6A19DD0691DA",
		INIT_0C => x"21EB3ED87BEC37D54472B0E5E25BF36545279038098D4DA358B490C8A190EA25",
		INIT_0D => x"D5EFDCD269B9BAE625D8A61B6D35C4EA3178CC7F033B844780CA21A8EA30F9E7",
		INIT_0E => x"0D7E5710C80A17AE3E94E7ADF8A8FC5248B1FEFBFAC66C71624609330E3E8904",
		INIT_0F => x"3C9B582201DCF6E595B28C0E8E215FAC49789D7AEC88D580B21C46F184CED1D3",
		INIT_10 => x"D5B42CDF726239F60D110304DAC9C61A56EE9A89751C6E2E0087CE8B7F4C7E30",
		INIT_11 => x"3057FA52E7A2F9449A7A558FAC2EAA6F4BA31B15E21A401C54C224CEEEBEF6C1",
		INIT_12 => x"BD66943F6FFF23FA20F0FC6F053AE56495CF3AD36744AF6C63AEDE5E10E77381",
		INIT_13 => x"EFC3093996D031C9A4BA92872052490DE752E982CF076C51233E94ADE6C79C48",
		INIT_14 => x"6A0E3332E0F48BE01C9681367E0112E4B1CD7CDF4A91F28092402F7911E00C00",
		INIT_15 => x"2065379A5480BE912A9CBBBAEA18820A6362DB186DBEF6259B3C4F130BDDF37E",
		INIT_16 => x"A46B44C3498C318496032F484BE2B9DC1259AB7BC8C8922A45F59D5BE06EDC2B",
		INIT_17 => x"DDB7994668E54D4C2C91077AFAEA1F82C4EA5F8FEFE42BAD830D05DAD46393CE",
		INIT_18 => x"EBED068DA6F64A2BF7CDE289101212B890C6D56AFEE0FA9FA2DC84036124DA1D",
		INIT_19 => x"936EF5307F7167F74A1AD431B6FBD9C01E7BD8D8AD36D9843385A1D7EEB571DF",
		INIT_1A => x"EBE6A8D98E0DA2CDB06BBF3B53F3C89E20CC1C7F8397C688B74D5CB93F7151B5",
		INIT_1B => x"35D5F68344AD2B6245D673BEFB95EC82F331016E9053BD44638378898E1A6350",
		INIT_1C => x"81C639129DD843C1CB954DFB02984B6D7C58EC808BBADD3FCC4F294D4F56617E",
		INIT_1D => x"FA5FF5EBDCBA56D7F73EA97B92D2DD519E624946A1FE2ACDCBE6C7F105816D3C",
		INIT_1E => x"33295926BB9FC23821BA08117AB9AD5BDA3EFED27C7179A5E44AC2653083C717",
		INIT_1F => x"7452E9E6EF10D35D9857D5B85957A73FEC8F1F1D1895EFDA181476AA4BF7BCAC",
		INIT_20 => x"5FCC2636863DAE1AE74B0200384734ED5B85063906D76A40FE1FE0B140A26059",
		INIT_21 => x"FC5BAC01FA4D9A9B4EBC5EECC940C45EA0AF8FC81D5D7F393B04A77D1D6C01BF",
		INIT_22 => x"0B93A9C098EBE8FB7331697B52C99E97118F751F0D5F28140D737F13C8689C73",
		INIT_23 => x"9C738545364BE19FBC383D6B8D71550A423EF0B178F4969921E6B4C91EF546C3",
		INIT_24 => x"966F49583E447287B4BB0C42EB753F515925AB27D21E1FB4F0B62B8FB7A59D33",
		INIT_25 => x"DC73F3C9F3EE3E5121B5B14D5597961B62A28A0D1702E96558ED9BC034DDA1FF",
		INIT_26 => x"2C01E10921712A33480F86350E09B1C1A4ED00F570EE50C2D15AC539B92E23D6",
		INIT_27 => x"801C08D77F351B531C65C267DF23752F6C33262B50BE0A05454D20D864AE81F7",
		INIT_28 => x"78A7160CCF274115E4EFF611F80E7BB2C30555CABDC2954267307A9FAFF08C56",
		INIT_29 => x"76B9CBF5C0581F687A99F88CF54D542B3483E19129A422ABFD543EED6005013D",
		INIT_2A => x"685E87509429F292F329DC1AD5E33B1A6FAD5EA846C1630CE232FFEFB00A2B39",
		INIT_2B => x"0386445A97AB313F55B0DAE1B036082B23E4256EFECB12240FD3E50710982E6D",
		INIT_2C => x"CA00C277CDB82DE208CCD92B4663486541211BE7C23BD7959F5A6E74DDEB9ABE",
		INIT_2D => x"558BD8D9B0E250C1DA5E93B9097869C1EB8EBDFFCFD03E1F2D1C4EEE569BFA15",
		INIT_2E => x"F99A4AC22775C8FA82567F7419E8F1D383BD26A1D15063174CD406243EB0FC98",
		INIT_2F => x"3652D6464002122C94DB74BD76464E2CD274C9073925E97DFC6699247C997404",
		INIT_30 => x"45A2B5655FE1BC249095D0F560AAE00100F9FF0F9B756CDFD0073852AA1E8FB7",
		INIT_31 => x"9E2811DCD1B4AAEB572EC8CB992E47EDD22B54D07515647137092A7A069647F3",
		INIT_32 => x"CFC7EE31C7CADD0A76948306AE58C8F0EB631F52F9AD29CAE24105BB169EE3CF",
		INIT_33 => x"597B6E9EAB58C633C82D2A2436785413F2C5DB5FF817714E192086893F5BD274",
		INIT_34 => x"97FC0E7D446CB20985EC25D4278951978AC6F65C62288C11E914A6340234A21B",
		INIT_35 => x"4E392AC14E9FCDF4CF91335185C7CC2E3BA2DBE3295815308C7FF0A6C331FCE5",
		INIT_36 => x"CE1D8BC474C6789CC2D084895657C2C1087B1C8C101154B323FF259C42ECE555",
		INIT_37 => x"E9CAAF16E381F55DEF70DE1CA448EDFDC295D6ACCC4A52B988D2008BDD1A6F78",
		INIT_38 => x"BFFDEA297E388F60C4F0CA1BB5F5D25560917264A4A51D210AB9E86CEB20992B",
		INIT_39 => x"32A1563A918236CF32E8B3AA7DBE924BA2A208A92036A17013AB7F9A16F90555",
		INIT_3A => x"A61A983DF3242984BF5B928F2A01DEE653B491D57941B50BE005F04A4F84A095",
		INIT_3B => x"9B3D34D1874EC6E70C53C2ACB6FB923335A5D72F4BED08917E9E835AC3E106F3",
		INIT_3C => x"DC10073B1B3A3D2D90EC9CE7605BB430CAD9800236FAD90F0721F7DC93B4C4AB",
		INIT_3D => x"A8E55DF4D14EF4687F6A39D0D546B23BEC95DFC496F1DD4599002359D765D14E",
		INIT_3E => x"9090B4F607520D260A78FD5A00BE175FEE4842EB3DBBFE531F672C98BE355DB3",
		INIT_3F => x"1C428ED2CAF9B26D01CCE16B4D0FEC8E0F7213C51291C6E8085BA057921EBD39"
	)port map (
		DO   => doutout,			-- Port 16-bit Data Output
		DOP  => open,				-- Port 2-bit Parity Output
		ADDR => addrin,				-- Port 10-bit Address Input
		CLK  => clkin, 				-- Port Clock
		DI   => (others => '0'),	-- Port 16-bit Data Input
		DIP  => (others => '0'),	-- Port 2-bit parity Input
		EN   => '1',				-- Port RAM Enable Input
		SSR  => '0',				-- Port Synchronous Set/Reset Input
		WE   => '0'					-- Port Write Enable Input
	);
	-- End of FRAME0000_RAMB01 instantiation

end FRAME0000_A1;