--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
--	Grupo de Apoio ao Projeto de Hardware  - GAPH
--	Projeto X10GiGA - FINEP/PUCRS/TERACOM
--
--	M�dulo:	Mem�ria - Gerador de Frames - Prototipa��o
--	Autor:	Jeferson Camargo de Oliveira
--
-- 	FRAME:	0004
-- 	RAMB:	01
-- 	CONJ:	A
--
--	M�dulo gerado em 17 de July de 2008 �s 16h55min pelo
--	programa gerador de frames OTN do projeto X10GiGA.
--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

----Pragma translate_off
library unisim ;
use unisim.vcomponents.all ;
----Pragma translate_on

entity FRAME0004_A1 is
port(
		addr	: in  std_logic_vector(9 downto 0);	-- Barramento de endere�os da porta
		clk		: in  std_logic;					-- Entrada de clock para a porta
		dout	: out std_logic_vector(15 downto 0)	-- Sa�da de dados da porta
	);
end FRAME0004_A1;

architecture FRAME0004_A1 of FRAME0004_A1 is

	signal addrin	: std_logic_vector(9 downto 0);
	signal clkin	: std_logic;
	signal doutout	: std_logic_vector(15 downto 0);

	component RAMB16_S18 is
	generic(
		WRITE_MODE : string;
		INIT_00,INIT_01,INIT_02,INIT_03,INIT_04,INIT_05,INIT_06,INIT_07,
		INIT_08,INIT_09,INIT_0A,INIT_0B,INIT_0C,INIT_0D,INIT_0E,INIT_0F,
		INIT_10,INIT_11,INIT_12,INIT_13,INIT_14,INIT_15,INIT_16,INIT_17,
		INIT_18,INIT_19,INIT_1A,INIT_1B,INIT_1C,INIT_1D,INIT_1E,INIT_1F,
		INIT_20,INIT_21,INIT_22,INIT_23,INIT_24,INIT_25,INIT_26,INIT_27,
		INIT_28,INIT_29,INIT_2A,INIT_2B,INIT_2C,INIT_2D,INIT_2E,INIT_2F,
		INIT_30,INIT_31,INIT_32,INIT_33,INIT_34,INIT_35,INIT_36,INIT_37,
		INIT_38,INIT_39,INIT_3A,INIT_3B,INIT_3C,INIT_3D,INIT_3E,INIT_3F : bit_vector
	);
	port(
		DO   : out std_logic_vector(15 downto 0);	-- Port 16-bit Data Output
		DOP  : out std_logic_vector(1  downto 0);	-- Port 2-bit Parity Output
		ADDR : in  std_logic_vector(9  downto 0); 	-- Port 10-bit Address Input
		CLK  : in  std_logic;			 			-- Port Clock
		DI   : in  std_logic_vector(15 downto 0); 	-- Port 16-bit Data Input
		DIP  : in  std_logic_vector(1  downto 0); 	-- Port 2-bit parity Input
		EN   : in  std_logic;			 			-- Port RAM Enable Input
		SSR  : in  std_logic;			 			-- Port Synchronous Set/Reset Input
		WE   : in  std_logic			 			-- Port Write Enable Input
	);
	end component;

begin

	addrin <= addr;
	clkin  <= clk;
	dout   <= doutout;

	-- FRAME0004_RAMB01 instantiation
	FRAME0004_RAMB01 : RAMB16_S18
	generic map (

		-- The following generics are only necessary if you wish to change the default behavior.
		WRITE_MODE => "NO_CHANGE", 	-- WRITE_FIRST, READ_FIRST or NO_CHANGE

		-- The following generic INIT_xx declarations are only necessary
		-- if you wish to change the initial contents of the RAM to anything
		-- other than all zero's.
		INIT_00 => x"9FF4B15F733C5FF1141E19F73BBD4BA4EE394885AEAB2CB045A9715105D2F628",
		INIT_01 => x"69229DCA5AE6C2DEE33812DE753710287F29F62BEE1FCC78FFD8E5FB5139892D",
		INIT_02 => x"999870CEE1039A353FEF11436639FEBB73E5E2F1F390E03A6083D3A5BC3AD372",
		INIT_03 => x"03D47686B890401A5CC7A157E7DE9B4177E0DA3D08B5B3D6F45DD036468BB732",
		INIT_04 => x"B8339A76B7CAE4C6E05D1B9DFAD2B3B75A5B2086F36EE4F665F6C85830772C84",
		INIT_05 => x"54C7CEF9529D9FA1BAB4A9FABDF549D17A9CE0B4B5A4CFFD90030D86371BAEB1",
		INIT_06 => x"E9FA485F135E53A173FC87A3734F5F3DBBA827687390187C6EC0A8936F2A45E7",
		INIT_07 => x"30B5D5C69E8FDBF5B699FAA5BF0ACFD9E0F2E0A4C55697DEEB733BB6E2C9115D",
		INIT_08 => x"068DEB307A132737ABBC035230ACC36FAE6D01BC387D840EB5484E52FC11672C",
		INIT_09 => x"0E32E587280F088E885A3076EF3359FA1ECB55817C6EA968668F875DFA88C23F",
		INIT_0A => x"FF9DDE137110E7BFCB5A31E0EAD7BEBA565D397737520C398017F2C6F49A2463",
		INIT_0B => x"1D559309FD77241E9CD49D5EDBE8D690399BAB3B593C06194E57CBA72899F869",
		INIT_0C => x"0EE2E52B8F97366DE376B8600EDCBF0EA454605B720134DCFC4FE7510B92370E",
		INIT_0D => x"CDD0C0753CA869B60BB6A38BC748781381F876A3FAB5C5848B481A5DA0B39A81",
		INIT_0E => x"F45CCB0BDFA5551311D0D37BD58474426988711266D19BDC128E63BA158D39BA",
		INIT_0F => x"A8BB43010047C44D71B1BDBE3BBB824C8D2524381BB6E2D681D4DEC0819161EC",
		INIT_10 => x"3329C2A8A8982EADB7B27978E5BA94F2E6891DC2909A3F22B6B9A9CACE6080FE",
		INIT_11 => x"8855B2609558878B59C60C5258F03E491530FF2C6A74F5FC7AEAA6EE54C082F9",
		INIT_12 => x"4DC67847F50E67945C620D608CE201E049873C6ADAC99028D3625ABCFDD621CB",
		INIT_13 => x"D6A6134999F7CC73C5697274CE7821020E083857715F00D91BD5DD707CF182EB",
		INIT_14 => x"38D0C7E96AF2898318F44B09A62FB891217427375545AF27A76A043B0356928B",
		INIT_15 => x"E65736CCFD81EDB0F05E836B8F3055159A5BA532745D93D975BE7B8984055A8E",
		INIT_16 => x"2949BC3CA7AAFBE96159604C6033E8A2514C4CEA66A4E41F354A70A59A1D5C07",
		INIT_17 => x"778563B182B15A686E78A872D5C245D95CC3DCD1FAD20A62D5ED60BAC1D61260",
		INIT_18 => x"8E2DCE2D1B42BA373AF5EED541E88C4688701289256E53ED3FE9167C7B7C068C",
		INIT_19 => x"7B77E971A4736757A5170B764DBFBA2070CF63B6A4721139AF4686213179CA4D",
		INIT_1A => x"7547E0614D37832971D2E2162B0B88F8BDBF2D299C6F748B5DC210D1EB881D36",
		INIT_1B => x"F4A160728241A6AB137057713C69D0890119C4A65AFE61A0DAFBFA25F0403E37",
		INIT_1C => x"2FB042109201DCE18DC26CDDB6EE7E942403BC62A5C29DF97B811A1D0A8C8ADA",
		INIT_1D => x"263C0E82BAEED67FB0F3CDEB2274D85A256CE61EC4177961C767568D05B9561A",
		INIT_1E => x"86B3410985F981CBE7ED5EDCC4DE0470306AD3FCDC96FF3C8802E21839DBC354",
		INIT_1F => x"7452E9E6D4B5BDDA2E8B68638949E70775CD1FCB394C05E9ACEAB5A208C64FA8",
		INIT_20 => x"A66E9D5FFFA394A1EE20EDE1B0D637993F23415A5DD4D48253EEAD70DBED761F",
		INIT_21 => x"CE57752BDB53D37198F45953A38BEE962A4B8BE1D0AD0A83E47972CD67DA1925",
		INIT_22 => x"8FA9E9908C0218F859CED8FA1135418A3614965C4EF8200358CC19374D5A0428",
		INIT_23 => x"6E1A75627400D7F523117A3DF767AEDE4058BAF8AF729EE0C730AAA9A294F2DD",
		INIT_24 => x"E68619B2F2BD0C4BECD0B122C590FB28681B192C668D42082D5207C51577B697",
		INIT_25 => x"C90737BDF74340C5FB17C18C3052C328AD7E5494D6E749815AC3841C0CBEE9C2",
		INIT_26 => x"D2C3A4FE38083E271553A12BC025129874816FB72663450B324E2B23E44FE44D",
		INIT_27 => x"D6BD496D26CD8C725ED5672FDDEFCA04636795D55CB18AEED9EE247F418DD51F",
		INIT_28 => x"B7E057678D998B8F90047F0558999687B0F0358D19E99F389DFE13D2AD92BC23",
		INIT_29 => x"7E4E2224CAC0D4242EB45D4A641BF780509CF14EC0C66981CC746D7F33ED1DB1",
		INIT_2A => x"16959CA7060F06AFEBB2EBBC6A8B86C30D93B45683C3342F73E3BEC945B919FB",
		INIT_2B => x"2472209AAD7990C0395EB0ECC826B99F7D04C3C6C9867B04914DB4AC90933E68",
		INIT_2C => x"2A616BA54871E35498F78B0D510806715BBAD82B56F918D11A352D571BD5616E",
		INIT_2D => x"AC0FD5B3099751FC60DD7376F2F7576F75D69FC5362E2A415DBBD9341C64FAAE",
		INIT_2E => x"37DD7C7F2D3D61F4902F691A92EE9B2E0D92B6BA6BECDB1CE868DFB011F96D67",
		INIT_2F => x"0124582DB21D324D1C66FC3FCC4180A73DEF9FCD2C0A5201ECCD899F1E22CDA9",
		INIT_30 => x"EA48BC6A76CC68AE38FF97DCCB6003B6910217BAE4746E8A761FE3BEA387D73F",
		INIT_31 => x"FAAE59FF9EF59F46F43EA034E59C50B9000145046169B17AB0306C80F799D52B",
		INIT_32 => x"AB4E197499A56E9D76B4D3667E493EB9373D493627534AB60CCEB45857E2BD39",
		INIT_33 => x"02A1D1D978891051B36CA7172AD2628ACA847A8FC6B4E33081320207D452F927",
		INIT_34 => x"0FBEEB22B3F3A735D3FC3BA39A58F1F4CCE740EAED55365A2864B3DED2C35610",
		INIT_35 => x"6D2912A16708D8BE793FD784E5CA0BF5C7FB0F0408605303FEC4E239A0F0C045",
		INIT_36 => x"1682D0A3159EA7048A2D5A98F569EDCBC7CEB532A332515FCB83844BFC62FDDA",
		INIT_37 => x"4AD85A76E8B69E368104AB6C25307E9A8061B658E43C55D6AC4D92EF225A17C8",
		INIT_38 => x"1ADF1E4F944D1E80B20D35F1CCBFC3E7E2D41F1D9AF66D1C68822C2A575AA5F2",
		INIT_39 => x"47F4F585BD953DE5DC6250594EBB1A826667F6643F7821EDC86284441B7FBEED",
		INIT_3A => x"2DD8FAF8B22604E4391310C9EFF9EF7C9952C67291A4E76E30E970FF54999991",
		INIT_3B => x"9D92DFB3C38827723454D216879D77BDB7705D85ABC2943BD97B4D31CBDC8FBB",
		INIT_3C => x"F83517056291A8D282B38634D8EED7826786B282AAB14065691E03DCC37894CE",
		INIT_3D => x"DF7E9DDE3EF925AEF29D5411EBD5C8A3E148559B91563DFCF18C7BAA7DEBF516",
		INIT_3E => x"476E0B7D6862643D6B4FCC178D5D8B7FAF389A6FF80F0D9D5B50D174D7C790E3",
		INIT_3F => x"7C0B9250CAF9B26D04132CC225686FCE5A80DC3FFBADEB43577F3272AF283EB0"
	)port map (
		DO   => doutout,			-- Port 16-bit Data Output
		DOP  => open,				-- Port 2-bit Parity Output
		ADDR => addrin,				-- Port 10-bit Address Input
		CLK  => clkin, 				-- Port Clock
		DI   => (others => '0'),	-- Port 16-bit Data Input
		DIP  => (others => '0'),	-- Port 2-bit parity Input
		EN   => '1',				-- Port RAM Enable Input
		SSR  => '0',				-- Port Synchronous Set/Reset Input
		WE   => '0'					-- Port Write Enable Input
	);
	-- End of FRAME0004_RAMB01 instantiation

end FRAME0004_A1;