--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
--	Grupo de Apoio ao Projeto de Hardware  - GAPH
--	Projeto X10GiGA - FINEP/PUCRS/TERACOM
--
--	M�dulo:	Mem�ria - Gerador de Frames - Prototipa��o
--	Autor:	Jeferson Camargo de Oliveira
--
-- 	FRAME:	0003
-- 	RAMB:	00
-- 	CONJ:	A
--
--	M�dulo gerado em 17 de July de 2008 �s 16h55min pelo
--	programa gerador de frames OTN do projeto X10GiGA.
--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

----Pragma translate_off
library unisim ;
use unisim.vcomponents.all ;
----Pragma translate_on

entity FRAME0003_A0 is
port(
		addr	: in  std_logic_vector(9 downto 0);	-- Barramento de endere�os da porta
		clk		: in  std_logic;					-- Entrada de clock para a porta
		dout	: out std_logic_vector(15 downto 0)	-- Sa�da de dados da porta
	);
end FRAME0003_A0;

architecture FRAME0003_A0 of FRAME0003_A0 is

	signal addrin	: std_logic_vector(9 downto 0);
	signal clkin	: std_logic;
	signal doutout	: std_logic_vector(15 downto 0);

	component RAMB16_S18 is
	generic(
		WRITE_MODE : string;
		INIT_00,INIT_01,INIT_02,INIT_03,INIT_04,INIT_05,INIT_06,INIT_07,
		INIT_08,INIT_09,INIT_0A,INIT_0B,INIT_0C,INIT_0D,INIT_0E,INIT_0F,
		INIT_10,INIT_11,INIT_12,INIT_13,INIT_14,INIT_15,INIT_16,INIT_17,
		INIT_18,INIT_19,INIT_1A,INIT_1B,INIT_1C,INIT_1D,INIT_1E,INIT_1F,
		INIT_20,INIT_21,INIT_22,INIT_23,INIT_24,INIT_25,INIT_26,INIT_27,
		INIT_28,INIT_29,INIT_2A,INIT_2B,INIT_2C,INIT_2D,INIT_2E,INIT_2F,
		INIT_30,INIT_31,INIT_32,INIT_33,INIT_34,INIT_35,INIT_36,INIT_37,
		INIT_38,INIT_39,INIT_3A,INIT_3B,INIT_3C,INIT_3D,INIT_3E,INIT_3F : bit_vector
	);
	port(
		DO   : out std_logic_vector(15 downto 0);	-- Port 16-bit Data Output
		DOP  : out std_logic_vector(1  downto 0);	-- Port 2-bit Parity Output
		ADDR : in  std_logic_vector(9  downto 0); 	-- Port 10-bit Address Input
		CLK  : in  std_logic;			 			-- Port Clock
		DI   : in  std_logic_vector(15 downto 0); 	-- Port 16-bit Data Input
		DIP  : in  std_logic_vector(1  downto 0); 	-- Port 2-bit parity Input
		EN   : in  std_logic;			 			-- Port RAM Enable Input
		SSR  : in  std_logic;			 			-- Port Synchronous Set/Reset Input
		WE   : in  std_logic			 			-- Port Write Enable Input
	);
	end component;

begin

	addrin <= addr;
	clkin  <= clk;
	dout   <= doutout;

	-- FRAME0003_RAMB00 instantiation
	FRAME0003_RAMB00 : RAMB16_S18
	generic map (

		-- The following generics are only necessary if you wish to change the default behavior.
		WRITE_MODE => "NO_CHANGE", 	-- WRITE_FIRST, READ_FIRST or NO_CHANGE

		-- The following generic INIT_xx declarations are only necessary
		-- if you wish to change the initial contents of the RAM to anything
		-- other than all zero's.
		INIT_00 => x"C854A34B328DB1A5A0FAD92E58F8A7BD3DBABFF17AAF45A9A0057A8B4E91F6F6",
		INIT_01 => x"1B7564BB8242F9CF73087824F408C77D3E6C8224011BB1350B16C1DD6B2F68C5",
		INIT_02 => x"6E9C8BDE8312F1329F8B46FB3AB12080DFC7248304EFB77B552A9DD41537194C",
		INIT_03 => x"6DAB81B24CA3B87F21D74E8B3B76AA165A3A12B08824F90A42CAF221DB1B2795",
		INIT_04 => x"011D9B49F2016ABBD13204043C325F7D3D96EA5A4F4D1F3E566BEE058F8B4112",
		INIT_05 => x"9E025E0B480A732C141B12DFAB1BA5B545D199E07402392A667A1C37CB457D12",
		INIT_06 => x"C1EDC87411E82E0E01259BB80BD5C6A6BF5EED0498CB6091716AD22B550F794E",
		INIT_07 => x"F1206BFDEF0E0B2969F17DB1ADB8B64B2A98FB93A3E09979DD9C5B5982842045",
		INIT_08 => x"7BD4D6A991D80BB9BF9314FA2E883036C918FC8C64BDF2A398D03A6D668DD200",
		INIT_09 => x"DCAA7B68EA29A2CC54CB409FD8DCE6AF2D050C5DA2AA0998767038372D1F0198",
		INIT_0A => x"2E0B680A2145D3164F765A92028F7F45E3F9630F79F826140232C80356790DD7",
		INIT_0B => x"EFD960B89B37A66B46ECA2988603FA011492302CF191A8110EF324D12EF3650B",
		INIT_0C => x"A67185655C8545600A535D91B519C956A6C228C77E087287E5064F9F0E5BF056",
		INIT_0D => x"80428AFA9DE9C73B3B7FC4C58FBB1DD30EAA647F7C67E8C8AFCB7A91C6CE7F6B",
		INIT_0E => x"C7B381BE4E4B8E8E39A64F793C225BF8B5FBBEA4065D6C056E15B2A342E1ABAE",
		INIT_0F => x"B17FA209EFD7ED34C30D8AC74C77171AF14D6D550CC0C12287CD86990149D43A",
		INIT_10 => x"1B71ED1B13C073DC6C3E8A7D1B665B26CC40D3D94ABE1A6FC768F76A5190D055",
		INIT_11 => x"A4E8B63266ED1037C6F0E7E614B752C81EFEF5CED5104FF06C22BC3A222B2573",
		INIT_12 => x"1F3329E43518334F7FFB9B5BB439341F530F8293BD4174CEE3B8F9154C07EBAC",
		INIT_13 => x"131A16E23501AECE2662D36F91B1594B34883CF029D93EB5EF1B9993A2474ACC",
		INIT_14 => x"B96C701F3609B39AF6EB74CA024E47F23FABDA3D200143A6DB93E958F2B4F178",
		INIT_15 => x"B3E6AE318C493E8E10BA2EA83CA7E540F08518B86CC72F9A8C80B6E7CBA684A4",
		INIT_16 => x"1517E9D5D345C486138FAD7FC0BDC1980368E838681356151015DE3A94E36582",
		INIT_17 => x"560F312348E309BD1C59D60788B79058918E277E44C676B414D71C5154F32301",
		INIT_18 => x"8551875CEA269C0E3DF999471099910AC7FEB71160F88D07801F0D4F59FDB123",
		INIT_19 => x"D9258B57F7192F845399A272AB778C9E4764FCDE5C14CDEB507F6C15A806C247",
		INIT_1A => x"1BE2FE78151AAD00EC8DD392DDCEA1F75E39BA515ED087E31B234F5BEFC297BF",
		INIT_1B => x"522844445D1E501D2D5787B18564711E1D84BAC18B6382237F1B8F981C25EFFF",
		INIT_1C => x"392316D1B92525FAD05F213899808637901F0A31780E0ED984FF71275C1E3A0B",
		INIT_1D => x"7F09D55C2EC4D0A3C7EE0C0FE23AA2B2A5D0ED7A33A039F52CD4CCD866E64B0B",
		INIT_1E => x"33455E851EAC0C2B2A35C09872AA2E83F60D0A4FA43057EEBDAA58B70D40844E",
		INIT_1F => x"E3C3B557B030121325F6768EE90BD5A18DB6318C4DA5266499A655BBD22C9195",
		INIT_20 => x"92823509A279134B4E89C02FD4AEE538554F1D43558D395D4A2B0A882CE6C2B1",
		INIT_21 => x"931563CA7A8AFED77F98CAE69034D33A2899C59C1405CF89151BC3948BFFD939",
		INIT_22 => x"20610EEDC7A7C1EE13818E318CA8C94FB162470E104B5FE89498BC6414733A51",
		INIT_23 => x"EE3830F4D9DD6AF2DE04D6698A61BB9D1F008BB45A5DE13D34165904F4ABBA9C",
		INIT_24 => x"57CBD5FBF12EF8AC2802D1D70B0EB3D378BADBB25CF1167214CAF03D8AA05AA6",
		INIT_25 => x"331361802DDF3C14B5EED3057B9FC144463EBA8C922CFE147BB4F45F34E428A7",
		INIT_26 => x"FC41518CC4B5E8F4893E6E7C8A7D7B54D1B0FFB9CF81A61FD14E74E4AC981D65",
		INIT_27 => x"3BA2985119856A0468B29B930168053C7025F8222D2526248F6F047642C081CC",
		INIT_28 => x"AC862D9320D3A4EC8591D041B92280A07D19DFA070B0E62B36B39909F1E8A73D",
		INIT_29 => x"14D79E3C119DBEFC9CC422AC2A4D47F14D91EA2AF29BBEB3F29A90FE0A2E3AD8",
		INIT_2A => x"BE6ACE5CE56989B8AFF9738BFC007E04F6F30CC421794D211B968E52F2FE57E9",
		INIT_2B => x"AA8B838C089513069D590F51EADBDDE4F2E2748E4C8792B66B5FEA1714E38D5B",
		INIT_2C => x"1DC736A0F0F88CA7ACACEBA09414627AF35282256323F2646959889E5DC81D32",
		INIT_2D => x"FC562C5C58D9EB17393355EB3EB8B1AD88641059E729F0AF7EF76D3ABD06DA4B",
		INIT_2E => x"11E6579342A1BF859AC2EEF98D79F27078D1EAFA2D8F7A8BFD4E110FE6405EFD",
		INIT_2F => x"341E7B5CF2DA3C5BC7F06F710A5A75C9E4189ABF0E2F8F3DF4D873A801B39F82",
		INIT_30 => x"F64D418F67602BBF2AD57CC02E91F5756761A3BEDFB3C923F0555E2C1923A137",
		INIT_31 => x"DD8E43FFA1997FED739C28FA075015B059A9EF75873811E728F198F928B74850",
		INIT_32 => x"EBE4C5875530DE4DA8C42BB9CF2A7C8BDE691D55B513D17D630546E560102CAE",
		INIT_33 => x"792428DF263C33C9AF62D79E51287A0B31F78C8DC3BFB22A3A6CB17A7EF63B36",
		INIT_34 => x"7F22CC48C9EF2ACA2A48F50DA5FBF603F4307A3F98A83BBACF863A0FB5C2494D",
		INIT_35 => x"45390DC643DBED9CA2A84E69FF02187F809E6AFCC664988AFFC9FB9C0C9E5F01",
		INIT_36 => x"CEF89B1DAC9E39ACA461005B1481BF5117FCB3A84086F7D0B0A2C7330A32CD22",
		INIT_37 => x"D1E205E89E3F2E361127C340FFA96CE21E11F5DD57DAF9724C8AA21D7A1C328D",
		INIT_38 => x"7CF545B4B7AD08C31A8D42C9E004D53FA378C7F46262C7995D58E034572593BB",
		INIT_39 => x"1A1DF61A67DBC7BB34C355810B1BE877911A4424C6821109EA816282CCF8403A",
		INIT_3A => x"CBC0251C5B72EE1389ED8BE2F8E8B6C535BD247540CB26B11BB25B73AC98ED08",
		INIT_3B => x"DC7251DA7460B6E8BCD0DD2472E1DA53C003CF5D648E780375C54D1AA53C38EE",
		INIT_3C => x"834AA961616CF65E0F0CC09ED8C68186E8240769D3BD64EDCF35A38C27C3F095",
		INIT_3D => x"7E658DD6D114C544F0613AC3497B1C47B97BE955273CD6EDAD10FBB4EF5C149E",
		INIT_3E => x"D375C70FD6DC0018E523C81A469F88FB7E7EAC024BC0194A025B6EF0D66E9EC9",
		INIT_3F => x"E5FDE8B9ADB671420E31E9856C0E84605A0DCD4B97CC9F2A6D6B04BB8441CA64"
	)port map (
		DO   => doutout,			-- Port 16-bit Data Output
		DOP  => open,				-- Port 2-bit Parity Output
		ADDR => addrin,				-- Port 10-bit Address Input
		CLK  => clkin, 				-- Port Clock
		DI   => (others => '0'),	-- Port 16-bit Data Input
		DIP  => (others => '0'),	-- Port 2-bit parity Input
		EN   => '1',				-- Port RAM Enable Input
		SSR  => '0',				-- Port Synchronous Set/Reset Input
		WE   => '0'					-- Port Write Enable Input
	);
	-- End of FRAME0003_RAMB00 instantiation

end FRAME0003_A0;