--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
--	Grupo de Apoio ao Projeto de Hardware  - GAPH
--	Projeto X10GiGA - FINEP/PUCRS/TERACOM
--
--	M�dulo:	Mem�ria - Gerador de Frames - Prototipa��o
--	Autor:	Jeferson Camargo de Oliveira
--
-- 	FRAME:	0004
-- 	RAMB:	02
-- 	CONJ:	B
--
--	M�dulo gerado em 17 de July de 2008 �s 16h55min pelo
--	programa gerador de frames OTN do projeto X10GiGA.
--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

----Pragma translate_off
library unisim ;
use unisim.vcomponents.all ;
----Pragma translate_on

entity FRAME0004_B2 is
port(
		addr	: in  std_logic_vector(9 downto 0);	-- Barramento de endere�os da porta
		clk		: in  std_logic;					-- Entrada de clock para a porta
		dout	: out std_logic_vector(15 downto 0)	-- Sa�da de dados da porta
	);
end FRAME0004_B2;

architecture FRAME0004_B2 of FRAME0004_B2 is

	signal addrin	: std_logic_vector(9 downto 0);
	signal clkin	: std_logic;
	signal doutout	: std_logic_vector(15 downto 0);

	component RAMB16_S18 is
	generic(
		WRITE_MODE : string;
		INIT_00,INIT_01,INIT_02,INIT_03,INIT_04,INIT_05,INIT_06,INIT_07,
		INIT_08,INIT_09,INIT_0A,INIT_0B,INIT_0C,INIT_0D,INIT_0E,INIT_0F,
		INIT_10,INIT_11,INIT_12,INIT_13,INIT_14,INIT_15,INIT_16,INIT_17,
		INIT_18,INIT_19,INIT_1A,INIT_1B,INIT_1C,INIT_1D,INIT_1E,INIT_1F,
		INIT_20,INIT_21,INIT_22,INIT_23,INIT_24,INIT_25,INIT_26,INIT_27,
		INIT_28,INIT_29,INIT_2A,INIT_2B,INIT_2C,INIT_2D,INIT_2E,INIT_2F,
		INIT_30,INIT_31,INIT_32,INIT_33,INIT_34,INIT_35,INIT_36,INIT_37,
		INIT_38,INIT_39,INIT_3A,INIT_3B,INIT_3C,INIT_3D,INIT_3E,INIT_3F : bit_vector
	);
	port(
		DO   : out std_logic_vector(15 downto 0);	-- Port 16-bit Data Output
		DOP  : out std_logic_vector(1  downto 0);	-- Port 2-bit Parity Output
		ADDR : in  std_logic_vector(9  downto 0); 	-- Port 10-bit Address Input
		CLK  : in  std_logic;			 			-- Port Clock
		DI   : in  std_logic_vector(15 downto 0); 	-- Port 16-bit Data Input
		DIP  : in  std_logic_vector(1  downto 0); 	-- Port 2-bit parity Input
		EN   : in  std_logic;			 			-- Port RAM Enable Input
		SSR  : in  std_logic;			 			-- Port Synchronous Set/Reset Input
		WE   : in  std_logic			 			-- Port Write Enable Input
	);
	end component;

begin

	addrin <= addr;
	clkin  <= clk;
	dout   <= doutout;

	-- FRAME0004_RAMB06 instantiation
	FRAME0004_RAMB06 : RAMB16_S18
	generic map (

		-- The following generics are only necessary if you wish to change the default behavior.
		WRITE_MODE => "NO_CHANGE", 	-- WRITE_FIRST, READ_FIRST or NO_CHANGE

		-- The following generic INIT_xx declarations are only necessary
		-- if you wish to change the initial contents of the RAM to anything
		-- other than all zero's.
		INIT_00 => x"EBE10DC646A82989B95A091FB12E48CE52CDDC399D1C2ED2A22082F86CF69ED5",
		INIT_01 => x"85FCD695AB5D290C68B394AC81C6D55245240EF0419C781C180EECAC52FB4352",
		INIT_02 => x"5E50A2F5402CC6DC7BBFA17DA3E81C18365EEEF28549BF8F6AE3ED6E5F24C9DC",
		INIT_03 => x"374D1466B0EB5CA8FC721B0DD07834B5438972BB79D5418124D299A55C14F3B9",
		INIT_04 => x"ACAAADF8C3E2F403651094EDBBAA5A77D9C7B5FC26AD36A06D8F29DAF5CAA092",
		INIT_05 => x"6DF82FEE42AFDCEBFC69F27F6D7EA180C520A8D5A04F7F8E8B450E326AE7F799",
		INIT_06 => x"5DD18856E4FFF5175FB26D4A2D766224E5E30FF92ABAD618A5DF19D5563C6661",
		INIT_07 => x"9F8B748F3C7E0B4C5A7B5A1A0013E9C195D74492AA11BCAF0CB7C27543B5AEE3",
		INIT_08 => x"DB336C8494EA15BD129CB9B35784607EF84EB6E55862AF616AB1D375F151EE70",
		INIT_09 => x"DDB752FF65F77C8F5470EC823BF18C9EE5440DD9561986032D4F0A549B661339",
		INIT_0A => x"0CD3AB004C5130D4E53BC31663D4A3C7DD172327F0AD79087C5855E1EC1594C6",
		INIT_0B => x"A271DF316DCD402673BDF146DA7F612E5651A843F256E01968C4B7B2511459D4",
		INIT_0C => x"CDAB866E4E049CA937A569963D285AAA779FBC21E9B28153EE97B7B7C6FF4F3F",
		INIT_0D => x"0C83DADE9863EFE3634A1E814044E200FA0DF67B873ACBCF3F990593E6E205A4",
		INIT_0E => x"3D1F03DA4ECEB9F101CE67617E66761B983EB30ECDA45099BA276530D074D8F4",
		INIT_0F => x"7DE734A3E6E8DAC5B0E61BBB6BD56CC5709C5FE72E31D54FBFC7AB738389A4FA",
		INIT_10 => x"A99847AB5B0C0BCACD6BCD3322AEDFD99C511CDDDD192C23CA37F7C6F6D3A2C7",
		INIT_11 => x"8E116822C26B6A7D4E6D2C3F0B069B628A736A3E836A4AC8E0E6B6212E85AEC3",
		INIT_12 => x"88D565D5CC2809FEDA64CAF66E621625B12913BA7D75082DFB94B75BEE6BFC45",
		INIT_13 => x"C903044441B2048A89E901D6C57FD666E76CB57CB4A0B2464555E913F71C453F",
		INIT_14 => x"685524964C6E7917B944D5925684D20A95114EAAA6563DF1F30C106988F12CDE",
		INIT_15 => x"AB5651D4FEFF2AF5AE15AEBE22DB707B4E094C9F7B01C90E147C08F0A54A5F4C",
		INIT_16 => x"4312328470D955F0E2AB96470415EB34D7DD79929D578A0E87EDDAA040B99E1A",
		INIT_17 => x"30EE1119AC33DD160C21B56F1ED1646F2EF4FCA7013CECC30B0B3ABFFA1D3CBE",
		INIT_18 => x"A6D30A262A66E8FE3D7B408D3A0DA30771F919C73EB60AFA91992B40B0230480",
		INIT_19 => x"C418EF1FB8EDD405B82D55F441CA83492F948A7CD1B8F23806CCB5372CB8A0B5",
		INIT_1A => x"3E7666A7B026CD79CD7A5E0991E14493289ADB1E0ECF5EA405805770EB71B1F3",
		INIT_1B => x"4DD3C7BF582CA2694DE08DB0DC5344898E96CDDB27D30D7579909E37480AE55B",
		INIT_1C => x"C4F8D09F2AA146CFC0721F6B9DC0163DB8D9DFF2C7AE4F472E97BD02E5F7F46F",
		INIT_1D => x"8F912E3C158214E802FD214CF05D853FAA64C802C783B2226C087B5014372ADE",
		INIT_1E => x"2CADF676B023E1BEA04C23A24BFE03BC4DE51E4548FE39A48A10BC5744BEE541",
		INIT_1F => x"D740BB244D37C0AA72BFB4EECED6DBF58B4CAC040B8F0AD2132E6773E33B4583",
		INIT_20 => x"B7D3A3F162348DE990F92D9CE4FE6F1EFED4BA052C66B5B43A4E8E666C76AF3D",
		INIT_21 => x"9AB4E6D566BE0633EB858CC8142F3F8DCC1563476BE2BA9EC3E09FBC342F4723",
		INIT_22 => x"52D0E79E6669289EA340A7AF5BA1160E152B399659F9BFFFA98303E179FABD35",
		INIT_23 => x"E110306327265D1AFA654F3DD009BA70E29863E585AABD03501E1CE0FA672850",
		INIT_24 => x"A484F3787F354CB5DE3FB65E732D32EED76722B8F3D178332328B7BD4055B338",
		INIT_25 => x"E8136AB40B7DEA0CDC37B37BCD2000DFB92BF6C01E85BD323F1FBC786947A1E1",
		INIT_26 => x"3F799A5CEDF5755F88B2B9F5D20A031880391F5F48A889046258BDD5BE89F37B",
		INIT_27 => x"FB9C5C9DE3D5973BC8C56621C4313F40FA5C8AF4FC0F7431FF6DF6351BEEFD7B",
		INIT_28 => x"42ECD39195EDAC004F261BA5F9A4F3DB25B10A09179BDBFEFBFD4D6CFC530D39",
		INIT_29 => x"B8BC03D3FE7CDDAFCDDF8795A78B246CEA113D214FBAEB230E8781453183F5EA",
		INIT_2A => x"A3FADDBB70F94AE018EA5B7FD955F6882BD841FAEF6EC74D206117930BA238BF",
		INIT_2B => x"8CFD90876360A89C01FD7CCC100EEEF69362066EF675B7AA63A35F057D4AD49A",
		INIT_2C => x"EA5A03597E63A22A760DF9EE8E367595D157597AA735B7D8004FFC32741CB1E5",
		INIT_2D => x"F32AE57238186230EFC299A9E902D07E3E9424EC4EF42E6E77BBA9DB5875D638",
		INIT_2E => x"BFE3B64848AEA63ADDB8C62115A95CD66E3BAB48E0E817AEB3F8E670D01BEAD2",
		INIT_2F => x"CF86C4B7C95D982BE2CDE6DB04D3BE50FDE32DD56B573594806A8E96BC47F335",
		INIT_30 => x"4B306695C2E9937BA7DAB97ECE12E55743511D1A393729317F1BD5ADB17CBB92",
		INIT_31 => x"668DD4E4D5E5003B083E270E728824CB8B771569AFFAFADCEC32E3463B218A4B",
		INIT_32 => x"2D0B1A8C5789FA9D3A5AD7C8B0EFFECF5D5D7057D0ADF21A43DD777A7A847836",
		INIT_33 => x"E9C328C5355D084651EA14E1659CAD9E20CAEE93701BE1188D12D171EDEC55CC",
		INIT_34 => x"8B0176CE22550C9AE76EE062AA9488A73367F365B66B0D42E79CCED5BE163947",
		INIT_35 => x"CC164D728CFD6057586C075F8C52C6D231C0940EAC4683277DF33BA97F641B1B",
		INIT_36 => x"09B13BC798D712FA95F2136A4B55236509C0FF27BAEA911BAF28283E465D3E21",
		INIT_37 => x"8DDA40DA594F077538431F0FF5D2E9CA359B704D73B1C0DCE1C549E5CE0BAE80",
		INIT_38 => x"0483537FC95DBD375CE61B94410EF266EA09FF3BEFCCF63685215FB994F9FC16",
		INIT_39 => x"EDF0387671E4699D8D6CF8EBCBFDE880EF8BBE8984D1D0A38E15D609BE3394B4",
		INIT_3A => x"2EA6A8787B3E7CD22FB2106361207D541B25F833D31CD8AE68A5454818FB5A63",
		INIT_3B => x"BA7AC270E2FC57EF27CCBB9079AE9E9786BAA347BE62B0ACE259D5B1AC364A9F",
		INIT_3C => x"F46D3F2C6C8141772BA7A1410226F7F5648429DE83C816A1BF459E704D0E58A7",
		INIT_3D => x"CAFD2746701C51606BD689E298AAF24E0AEF4179A3B9E625DE5B84E88DA121A7",
		INIT_3E => x"138A98E76A1DD3FA8C7426B0F938DF97297DDC9D115D31E96C237D25BD6278AB",
		INIT_3F => x"1111111111111111111111111111111131CE398538CFB28EB2DD1E3E4957CF1C"
	)port map (
		DO   => doutout,			-- Port 16-bit Data Output
		DOP  => open,				-- Port 2-bit Parity Output
		ADDR => addrin,				-- Port 10-bit Address Input
		CLK  => clkin, 				-- Port Clock
		DI   => (others => '0'),	-- Port 16-bit Data Input
		DIP  => (others => '0'),	-- Port 2-bit parity Input
		EN   => '1',				-- Port RAM Enable Input
		SSR  => '0',				-- Port Synchronous Set/Reset Input
		WE   => '0'					-- Port Write Enable Input
	);
	-- End of FRAME0004_RAMB06 instantiation

end FRAME0004_B2;