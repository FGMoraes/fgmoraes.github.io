--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
--	Grupo de Apoio ao Projeto de Hardware  - GAPH
--	Projeto X10GiGA - FINEP/PUCRS/TERACOM
--
--	M�dulo:	Mem�ria - Gerador de Frames - Prototipa��o
--	Autor:	Jeferson Camargo de Oliveira
--
-- 	FRAME:	0000
-- 	RAMB:	02
-- 	CONJ:	A
--
--	M�dulo gerado em 17 de July de 2008 �s 16h55min pelo
--	programa gerador de frames OTN do projeto X10GiGA.
--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

----Pragma translate_off
library unisim ;
use unisim.vcomponents.all ;
----Pragma translate_on

entity FRAME0000_A2 is
port(
		addr	: in  std_logic_vector(9 downto 0);	-- Barramento de endere�os da porta
		clk		: in  std_logic;					-- Entrada de clock para a porta
		dout	: out std_logic_vector(15 downto 0)	-- Sa�da de dados da porta
	);
end FRAME0000_A2;

architecture FRAME0000_A2 of FRAME0000_A2 is

	signal addrin	: std_logic_vector(9 downto 0);
	signal clkin	: std_logic;
	signal doutout	: std_logic_vector(15 downto 0);

	component RAMB16_S18 is
	generic(
		WRITE_MODE : string;
		INIT_00,INIT_01,INIT_02,INIT_03,INIT_04,INIT_05,INIT_06,INIT_07,
		INIT_08,INIT_09,INIT_0A,INIT_0B,INIT_0C,INIT_0D,INIT_0E,INIT_0F,
		INIT_10,INIT_11,INIT_12,INIT_13,INIT_14,INIT_15,INIT_16,INIT_17,
		INIT_18,INIT_19,INIT_1A,INIT_1B,INIT_1C,INIT_1D,INIT_1E,INIT_1F,
		INIT_20,INIT_21,INIT_22,INIT_23,INIT_24,INIT_25,INIT_26,INIT_27,
		INIT_28,INIT_29,INIT_2A,INIT_2B,INIT_2C,INIT_2D,INIT_2E,INIT_2F,
		INIT_30,INIT_31,INIT_32,INIT_33,INIT_34,INIT_35,INIT_36,INIT_37,
		INIT_38,INIT_39,INIT_3A,INIT_3B,INIT_3C,INIT_3D,INIT_3E,INIT_3F : bit_vector
	);
	port(
		DO   : out std_logic_vector(15 downto 0);	-- Port 16-bit Data Output
		DOP  : out std_logic_vector(1  downto 0);	-- Port 2-bit Parity Output
		ADDR : in  std_logic_vector(9  downto 0); 	-- Port 10-bit Address Input
		CLK  : in  std_logic;			 			-- Port Clock
		DI   : in  std_logic_vector(15 downto 0); 	-- Port 16-bit Data Input
		DIP  : in  std_logic_vector(1  downto 0); 	-- Port 2-bit parity Input
		EN   : in  std_logic;			 			-- Port RAM Enable Input
		SSR  : in  std_logic;			 			-- Port Synchronous Set/Reset Input
		WE   : in  std_logic			 			-- Port Write Enable Input
	);
	end component;

begin

	addrin <= addr;
	clkin  <= clk;
	dout   <= doutout;

	-- FRAME0000_RAMB02 instantiation
	FRAME0000_RAMB02 : RAMB16_S18
	generic map (

		-- The following generics are only necessary if you wish to change the default behavior.
		WRITE_MODE => "NO_CHANGE", 	-- WRITE_FIRST, READ_FIRST or NO_CHANGE

		-- The following generic INIT_xx declarations are only necessary
		-- if you wish to change the initial contents of the RAM to anything
		-- other than all zero's.
		INIT_00 => x"FFCE6EA5FCA99DFF89417A4505ADD3E83891008F0E6B54EBA8B23813131F2828",
		INIT_01 => x"57A154D860B458D0622794338E41563F13FBF4F1EE05F2DAD7C56430A4035FF7",
		INIT_02 => x"F91719BFD6AF01DE191A8C9C9555961A788A5AD7583210C0CE630AE02834CC6A",
		INIT_03 => x"DEC404E8B3C5A04206C0579C684E9EBFF99DEE4639B3E31D278D40F551875411",
		INIT_04 => x"9F84D11272F498ED8FCDE2823D5B346BE2558D3E973E4CC6730DA40C33B80633",
		INIT_05 => x"DFE7FCD6C6A01FDC0153783AE237C910B69D879C620CD9AF3774A3656D324FBE",
		INIT_06 => x"FFB74A954A038AEE8FC1BF378577B4B73DF59CB4021C06FDC626911F7DD5BC01",
		INIT_07 => x"1DAEC0C6C17404179B60D4EAE951ABE3C2E11FA30321550051546FD36DB89ED1",
		INIT_08 => x"5C571DD3E76499373F50D4B7C21244EC1A6906576703D4F0FBF7146EE923768F",
		INIT_09 => x"772325FD22C7998D4BDA097A746921A7733E67EEAC13891896F88837415904E2",
		INIT_0A => x"C35011F0691A7AA8B38B6ED1D22CDBD4E299C5B7F126ACEFFA3D7B0FAB7FF5F4",
		INIT_0B => x"96A2BCA5CF35F7AF192D5B9C0FD512F18BEEEFB4FE4B3A6DF21C9E4D259BD18D",
		INIT_0C => x"668FD70D8E3EE79A8C32E50CFC0185E20B45D103299577C0977FB3509C4C127E",
		INIT_0D => x"76A397ED379BB8AE8F498377C451BF8F9B93756F3A5FE0651BC1732487000776",
		INIT_0E => x"D4BC59C974C3A18C9A650B434255AF8F0EB9DEC8AAC7896AC22B45CEE8BE64FE",
		INIT_0F => x"EB4759BF808A9D8226F7E52DBBB96B072CF2B50C313F7567DE835C2E5CF110D9",
		INIT_10 => x"2FDF36C38FF32BB7B5C6460EFF3FDF720774A63418B8FEAD474DAA08F615FF5B",
		INIT_11 => x"E6AF19F061F00B04EA74E769818FD2FB5277AE1FA2671B1CC13E8C09CE6DA943",
		INIT_12 => x"80D752B8672E4A590BC33919256573CB86A6C9F7BC2166B3D51E8A641E73062E",
		INIT_13 => x"D09A2482BC9A7A074B535BFA0B38106D4CA5CD446E59DE635137DD813FCF183A",
		INIT_14 => x"5DFCDB2A39D7799D495BE5831FD6C0D0B1228AF7A03402770689C79E5153FF4F",
		INIT_15 => x"EB64E61F29B0C27FB7DE69E6871B4AB68EE3D83424F9A6E62946E1D056784357",
		INIT_16 => x"A4C021C96017955DA430C4ACA64FE0DDDF7A97D27FF12DDD1137290BB938ADEC",
		INIT_17 => x"64EC60137F8C9C8986F2800B073589641F775729382E623071ADB0E05113E390",
		INIT_18 => x"B55768CDD51765ACBA8BD88D3E3062ECA62A3043206810755F602A3C9CDC3C06",
		INIT_19 => x"8483473A4A1FEA80C1A074023A7038016BC7494B4F67BAB637903062BF87FAF2",
		INIT_1A => x"D4D6FDA514E44822FC78DA4B0CA30B52984C82327B42E5F4F54531AA9C23E976",
		INIT_1B => x"3FE87D34C62827023D37DFB529061A0B08498072C8F959342A19ED3375378C8C",
		INIT_1C => x"4C4CB2E1B20074CFE4E479CF2AE8938E304E37022FDC4301056C838F687F7329",
		INIT_1D => x"4D073042B0EFAD9B2F6C400D01CFB069853EC893701D59BCEF3DFBBE5DA0D7FB",
		INIT_1E => x"899F83B2DDD525904B9952B93C6167C94D704959FE67E6A9C49CB78FAF936D82",
		INIT_1F => x"DCB1CB430B576FFB64ED713A72048DA94A36E56D9070F191CDE1499D4F140019",
		INIT_20 => x"E23D6AA2295654B9CB0736E97ACFF9FF382F1A1909416544240849E9CF54145B",
		INIT_21 => x"61D865BB2E2CC26A848AF0C9E41B309382475C96AA5191612DFB55E7E343C153",
		INIT_22 => x"D758C7C412E3D4AE722FD2D57347ECDBC94FCECA5D6D0ACF2932949EC2947B9B",
		INIT_23 => x"A89A30E12CB2E0BD4345CFD0C8417A3C2797B55685EF0EEA4F27945E9CE79768",
		INIT_24 => x"4D9CDDE2148E1CD41DA4A0752A019F5604F04AD0F3D1838DB0D303AB443B5145",
		INIT_25 => x"775A9AB3B4A80B942964013EF216028D447ADC2948AF1B22AE6F686F01383E53",
		INIT_26 => x"3724F7E421F21F88E7F6A7B02535BBFD24312748DEFA621B28732596714BC2E2",
		INIT_27 => x"3A6503F63FF4C0B146B560B8A52DEB8AB221A4A75351D9AC460A58FB4DA6FB9B",
		INIT_28 => x"07BF743FE2BDE8169ADE46D9B76FC0195496BA34AF0FBA3B7CCF6B38D5F08C8A",
		INIT_29 => x"AE05F959DC87DC7981A29F81A4057F4CC78A26E8C90DF4D4DAD0597E2BB4F602",
		INIT_2A => x"8BC26BEBC5E2ADD6BCB094ADEF400E3A213D064156EE26461A4CF8F3995706F3",
		INIT_2B => x"9FB6EA2E638151E758F0822DAEF4C6E18DD0EBD3C2F47B00F6E63C9DA29A7B41",
		INIT_2C => x"56537220493A6076C0BF4F29618A05A0E8AD60E2265164CF110BFA37AF2ADA14",
		INIT_2D => x"0095641A37B10AC24A64DE1B45A09F351C5525FEEB45F7DE58F63AAC9C92D3C9",
		INIT_2E => x"A4411D7EA3FAEDE045E26C11CA6A5054BC01B01B0717CD63BD1751FC347E6139",
		INIT_2F => x"42004FC2EA6487BF2C656AAA62503590ADCCB818F40B10054913349EB50C8F04",
		INIT_30 => x"F3424E37153C7632856E38C1D54BF08500247F435D2D33C009605EAF539D8283",
		INIT_31 => x"C87AB0C745BC4F0AA6FC9F1428B4370E34C3ACAF9722AECC014A55778054DBE1",
		INIT_32 => x"BEA3B8DFA2CD694FB5D345C3F240976A68A462779EAAC87B07FDD9A740C7EF18",
		INIT_33 => x"BF1258D84D9D10D62D47672839E6AC0BD77E24AC15DA4F7CC10FBA889865315B",
		INIT_34 => x"732C5487BD36D25B6FE97755F54818A61B38DD511B654747A3D3773D50B800AA",
		INIT_35 => x"D5FB3758E073D861D7CB68385B759FCDFDD4DA2A319B5E325E734EE9E0B8212C",
		INIT_36 => x"3B1140FA592C7D95371E4B0221F3D0D661322B56F8445BD5A22034E66AC7E107",
		INIT_37 => x"E3D3846060916B0B2294649DC1554C697D8843EA71BCBC9C227FAB9877CE307F",
		INIT_38 => x"2F670B0A85EA21CC762FB773CFE280B737A2162A62AE864C167715F2CC00F3A2",
		INIT_39 => x"7848903DCB5A37B195D9CB4BCD2354ABB94259540E1C209536D42311EB7F9C6E",
		INIT_3A => x"90B810DC29C4C578D8D2937C8658777AB6DFC07E4B70EA91DAF6EDAEAFCC170D",
		INIT_3B => x"D9D245BC42B9484B7981F09BAA67004117DC4AA1C912AFEF7B2D1E5604979900",
		INIT_3C => x"092A751953606B74475E17175424B8DC67EB16304A7DA3E21E7BD93E6832557F",
		INIT_3D => x"3654899ED61EBC2BFC538DB571B1CEF60A1ADBE85DB6995D21ED59DC0D5C975C",
		INIT_3E => x"B713245ECADC9FDD3DB76637969FC60A0E59303A10C89C0AE10EA88B98C8A62F",
		INIT_3F => x"07DE8AA59BE9CF0F5CB2E77EB761FEB6984BCB4A631D85218D1E6BD9FB466B5D"
	)port map (
		DO   => doutout,			-- Port 16-bit Data Output
		DOP  => open,				-- Port 2-bit Parity Output
		ADDR => addrin,				-- Port 10-bit Address Input
		CLK  => clkin, 				-- Port Clock
		DI   => (others => '0'),	-- Port 16-bit Data Input
		DIP  => (others => '0'),	-- Port 2-bit parity Input
		EN   => '1',				-- Port RAM Enable Input
		SSR  => '0',				-- Port Synchronous Set/Reset Input
		WE   => '0'					-- Port Write Enable Input
	);
	-- End of FRAME0000_RAMB02 instantiation

end FRAME0000_A2;