--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
--	Grupo de Apoio ao Projeto de Hardware  - GAPH
--	Projeto X10GiGA - FINEP/PUCRS/TERACOM
--
--	M�dulo:	Mem�ria - Gerador de Frames - Prototipa��o
--	Autor:	Jeferson Camargo de Oliveira
--
-- 	FRAME:	0004
-- 	RAMB:	02
-- 	CONJ:	A
--
--	M�dulo gerado em 17 de July de 2008 �s 16h55min pelo
--	programa gerador de frames OTN do projeto X10GiGA.
--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

----Pragma translate_off
library unisim ;
use unisim.vcomponents.all ;
----Pragma translate_on

entity FRAME0004_A2 is
port(
		addr	: in  std_logic_vector(9 downto 0);	-- Barramento de endere�os da porta
		clk		: in  std_logic;					-- Entrada de clock para a porta
		dout	: out std_logic_vector(15 downto 0)	-- Sa�da de dados da porta
	);
end FRAME0004_A2;

architecture FRAME0004_A2 of FRAME0004_A2 is

	signal addrin	: std_logic_vector(9 downto 0);
	signal clkin	: std_logic;
	signal doutout	: std_logic_vector(15 downto 0);

	component RAMB16_S18 is
	generic(
		WRITE_MODE : string;
		INIT_00,INIT_01,INIT_02,INIT_03,INIT_04,INIT_05,INIT_06,INIT_07,
		INIT_08,INIT_09,INIT_0A,INIT_0B,INIT_0C,INIT_0D,INIT_0E,INIT_0F,
		INIT_10,INIT_11,INIT_12,INIT_13,INIT_14,INIT_15,INIT_16,INIT_17,
		INIT_18,INIT_19,INIT_1A,INIT_1B,INIT_1C,INIT_1D,INIT_1E,INIT_1F,
		INIT_20,INIT_21,INIT_22,INIT_23,INIT_24,INIT_25,INIT_26,INIT_27,
		INIT_28,INIT_29,INIT_2A,INIT_2B,INIT_2C,INIT_2D,INIT_2E,INIT_2F,
		INIT_30,INIT_31,INIT_32,INIT_33,INIT_34,INIT_35,INIT_36,INIT_37,
		INIT_38,INIT_39,INIT_3A,INIT_3B,INIT_3C,INIT_3D,INIT_3E,INIT_3F : bit_vector
	);
	port(
		DO   : out std_logic_vector(15 downto 0);	-- Port 16-bit Data Output
		DOP  : out std_logic_vector(1  downto 0);	-- Port 2-bit Parity Output
		ADDR : in  std_logic_vector(9  downto 0); 	-- Port 10-bit Address Input
		CLK  : in  std_logic;			 			-- Port Clock
		DI   : in  std_logic_vector(15 downto 0); 	-- Port 16-bit Data Input
		DIP  : in  std_logic_vector(1  downto 0); 	-- Port 2-bit parity Input
		EN   : in  std_logic;			 			-- Port RAM Enable Input
		SSR  : in  std_logic;			 			-- Port Synchronous Set/Reset Input
		WE   : in  std_logic			 			-- Port Write Enable Input
	);
	end component;

begin

	addrin <= addr;
	clkin  <= clk;
	dout   <= doutout;

	-- FRAME0004_RAMB02 instantiation
	FRAME0004_RAMB02 : RAMB16_S18
	generic map (

		-- The following generics are only necessary if you wish to change the default behavior.
		WRITE_MODE => "NO_CHANGE", 	-- WRITE_FIRST, READ_FIRST or NO_CHANGE

		-- The following generic INIT_xx declarations are only necessary
		-- if you wish to change the initial contents of the RAM to anything
		-- other than all zero's.
		INIT_00 => x"8EC9EF8DA600EA126F33D7E010CFC2C0C1814B18FD3F0226DDB47371131F2828",
		INIT_01 => x"03B63F1F3F547CB12FF8E986BA63FA58162C72D69F4FA6198F5FA57697E42763",
		INIT_02 => x"9F8D59D5DDCD309F587403BE09D904203225A97A62E74A509178F9E98F8A3751",
		INIT_03 => x"6010167188A766DA4EA642189063D11310923586A8BB2B87E023A82CDA71F9A2",
		INIT_04 => x"7619843995BEBF0F9C6598630399137EAE41F835797E557A0835BFB7E28B6207",
		INIT_05 => x"2413C8196D69028F47CE6B5987281D88A6C0BE27CD07F3AF3A1BB4EC017056F7",
		INIT_06 => x"1C11A36B049FFD123D98226A25B116914AE4A17C5CAC02A03F9D08B588C708E1",
		INIT_07 => x"F2033F0A91785750E6E96A1DD09A5EBAFB83BFBA7CCB8651429452A76E78BBDB",
		INIT_08 => x"2D6D53FA9C23F0BBA9CEBC846590F3296839BD6FACD54773A681E4EBB6FB388A",
		INIT_09 => x"0E694EB6029CDBB80898174E14962CDB1BE432C326CA7834003B43FDC0AA610E",
		INIT_0A => x"EEB79B92A0E6E3544D3D74BD0DF8A257A8857CE88D672A9115B9F804CF1133D7",
		INIT_0B => x"9762A3ACF4FC28242F8147D96782A575DBB75893A52A34B95168E1442B614132",
		INIT_0C => x"A693494EF4AFAD573937C788CA5E6A43FE5D05BD3207CCEE13E73DA038A857F4",
		INIT_0D => x"E744DD44E9609C1B9E39D2C728697393F4BD235874FFC96A9ACD9FBA21A6BAB4",
		INIT_0E => x"140C7F774C6B3549A903A2F46BFB6C85DFB78BE99EB4E2AEB9E76C7039318320",
		INIT_0F => x"5B8B4768E1DBA137E71AA1588D3D652C2328A23CA0FFB5DEAB487E0B786BC584",
		INIT_10 => x"3A106755D5366615CC83D3A5CFF9031A14683C09638D48EF95320FEF7C711883",
		INIT_11 => x"8DE5760C7B999F070BC7796B245A33B1448ACF99563A6FCE45EE96FD93FB5ABB",
		INIT_12 => x"1EA68060869C02C2006FC0C13D858595F3E4690C6B80082006585D2B2D560CDB",
		INIT_13 => x"2AFEB8801440BD028BBC63BB223AE7C23F84646DC4534B9A1C6C35D21DE568D7",
		INIT_14 => x"3B5F3401280C3625EC91DAC90DAF78B8A2A2B9BE15D8109750454B15BBD407F4",
		INIT_15 => x"8F743748644ABE9CABF4037C274D26561C2853B8EAD479A27743C726FDA2FF31",
		INIT_16 => x"D05FA4167C4F6DED7EA56F1C3734462B1D7B9ED3D90F7DC37A47D8431CAEF094",
		INIT_17 => x"64371D3766415DB414A056F9FDE377787AB79D8BF77F9EA556ECBA35720ED78D",
		INIT_18 => x"78022922AD1AE03C1891BD38173536F8718944D56844BF2233910340E8EA62EF",
		INIT_19 => x"9F601E363A664C6B16CD62F30E7C1DEC6A96583244EE7BA0A96DC6201F5837A2",
		INIT_1A => x"FC7C97BE3FFAF834699A4FC4660D0E0F4F07C8EB735F2E452E41DA473B5DA076",
		INIT_1B => x"8D2FCD413B4C11D8FCF35D96764BA67FB6A3C724A5A9520326BB96D00A0DD81A",
		INIT_1C => x"0E057B0B8F6AA9C680981F0E807BD99FD58FB58C165A733AA05CE71760AF8338",
		INIT_1D => x"FA5F24A43968EBB0A95D29A6C49B0A450D7716BF8BBB5EB16176D5F4F43AEE31",
		INIT_1E => x"E920A7AAA24F76F93E654989549EBE6D1801676A4537BD5588248F12FF665C68",
		INIT_1F => x"DCB1CB43E153274E1602E04E7221518C8B983B534F6715879859F10FF5534B9B",
		INIT_20 => x"5800477C39D8C5689699CE47473082582CE79D54BB08B3C62278B04E40B63B68",
		INIT_21 => x"2187B4220811781BDBE4C0345822A6C07EF2B23FC8F5C9013060A9A3CB8A7D61",
		INIT_22 => x"B367903EE05ED4646A6C2493A600BA284AAD8689ED3064AD98BFA2990198D80F",
		INIT_23 => x"64FB9DE32C673BFE3F3A9DBAE3CF9362D7725851CCFDB0DE6F77B941254B3628",
		INIT_24 => x"B9EEF088CE67489A31A72E0812AED84C17AAC3804644EF64C5CDC9FD75B9A9A0",
		INIT_25 => x"834138A571F6B7101834946110A603D3EE5E5C8F10AF3547FE5198FC09B9C555",
		INIT_26 => x"4C48851A9956E549C60CEF6A96D1B84D143E7ECD218EDFD6E7924686B0BDAE61",
		INIT_27 => x"6796107443F0897D55C2F0C97E6FDC372CE553E6720AD691FEEDBD484DE880FA",
		INIT_28 => x"AA10E0D295BAE3E933E3CBFDC0CA42CBBE39996C2C8ABBAC099A77C4CE4EE3B0",
		INIT_29 => x"311A7EF18570025C0E5BDC9D2EFD1C91389BF5C5526FFB856BC1C890C8BDF70D",
		INIT_2A => x"5628C3DBD281ED9363235CECC3DB04816A96300EDAF72A9602640C502BDE8919",
		INIT_2B => x"73961636A0BAAAFF14964FC666F2DDB0D1FFC26693BDBE4350E456DD06CD281E",
		INIT_2C => x"ACB1725BB9DB2D8987019CDEDEEEA65E4EC216E1D558423551A8B32DEB2D815E",
		INIT_2D => x"12B6DA15E25E69D10DDB65A32FF461794DFC10F19A44D351E50F9DEAC8AB6EB4",
		INIT_2E => x"6F81C38B98D0805521F31A15052D8371E83B4A3DDA72F9DB5B116E61D8DCD309",
		INIT_2F => x"32AACC0EFC8E117BCA8CD8D7B2F1056768034899273498542F7388F31558756C",
		INIT_30 => x"1AB8B9839ACFC4EDFF6074749A2D95E43B3FA9745CFF169A16832F6F26EDB54B",
		INIT_31 => x"F777153BA110CECA4E063FCDD53047B6098633525F19DF9C54997A0BAB1F19C5",
		INIT_32 => x"7B63DAAE9D5ACA4148BD49690E419893A209AC9995BFB59C86F58F101B0B3523",
		INIT_33 => x"7FF8030B31D02D7D0320101C09C3D4E34994CD351B8FAB57E558C4AE9AD97737",
		INIT_34 => x"B95300EF35077CFC33C2247D76E00AA1E7FF4B536E489F2B9D0C0DB22A2A97FE",
		INIT_35 => x"13D1FF167C4EC99233ADFABC12B828FB039D29F44988BA7D0763E4C3D61D7323",
		INIT_36 => x"FF438F19D71BF9A3253E8CE4141911D8292E467C927E0D62795BE53A951D7037",
		INIT_37 => x"DD999049EDC7108DFBAD8473D89BB580F83D5546AAC6C10286990FFEA27E5D92",
		INIT_38 => x"E3C8F1641046863290844E31591720B55C75A7F9FE95C90E70EAD7A5F6EE001D",
		INIT_39 => x"6D43ACC5181CA061F75778616CCAEB7B3A1EC1A04C40F50A313F5BAA86F5EA87",
		INIT_3A => x"DB0917D0B67EB1DFDEC70067C50033C2DA3432972A444BE3BE1F283DCAA14557",
		INIT_3B => x"6F4B3B657E36CA252090D460D2F1E0A8FC5F818023D2C7823D9775F287300847",
		INIT_3C => x"2B91A231212DB00896C8095D87FB8AD41C1D696A632282C91E86B370EEE9B21F",
		INIT_3D => x"8D1E68D226FB4FDF62BB33D44609A0B6A967817F795EB84802804A186A2B28E1",
		INIT_3E => x"578D7F6794FD427DF33F105BDDEF3E3165071C6EB62C27793AFAF4C8167A289D",
		INIT_3F => x"272E89489BE9CF0FF2707324C9B15FF49CA127288B494905CA38BF96CBDBECB9"
	)port map (
		DO   => doutout,			-- Port 16-bit Data Output
		DOP  => open,				-- Port 2-bit Parity Output
		ADDR => addrin,				-- Port 10-bit Address Input
		CLK  => clkin, 				-- Port Clock
		DI   => (others => '0'),	-- Port 16-bit Data Input
		DIP  => (others => '0'),	-- Port 2-bit parity Input
		EN   => '1',				-- Port RAM Enable Input
		SSR  => '0',				-- Port Synchronous Set/Reset Input
		WE   => '0'					-- Port Write Enable Input
	);
	-- End of FRAME0004_RAMB02 instantiation

end FRAME0004_A2;