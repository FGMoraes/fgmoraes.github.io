--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
--	Grupo de Apoio ao Projeto de Hardware  - GAPH
--	Projeto X10GiGA - FINEP/PUCRS/TERACOM
--
--	M�dulo:	Mem�ria - Gerador de Frames - Prototipa��o
--	Autor:	Jeferson Camargo de Oliveira
--
-- 	FRAME:	0002
-- 	RAMB:	02
-- 	CONJ:	B
--
--	M�dulo gerado em 17 de July de 2008 �s 16h55min pelo
--	programa gerador de frames OTN do projeto X10GiGA.
--++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

----Pragma translate_off
library unisim ;
use unisim.vcomponents.all ;
----Pragma translate_on

entity FRAME0002_B2 is
port(
		addr	: in  std_logic_vector(9 downto 0);	-- Barramento de endere�os da porta
		clk		: in  std_logic;					-- Entrada de clock para a porta
		dout	: out std_logic_vector(15 downto 0)	-- Sa�da de dados da porta
	);
end FRAME0002_B2;

architecture FRAME0002_B2 of FRAME0002_B2 is

	signal addrin	: std_logic_vector(9 downto 0);
	signal clkin	: std_logic;
	signal doutout	: std_logic_vector(15 downto 0);

	component RAMB16_S18 is
	generic(
		WRITE_MODE : string;
		INIT_00,INIT_01,INIT_02,INIT_03,INIT_04,INIT_05,INIT_06,INIT_07,
		INIT_08,INIT_09,INIT_0A,INIT_0B,INIT_0C,INIT_0D,INIT_0E,INIT_0F,
		INIT_10,INIT_11,INIT_12,INIT_13,INIT_14,INIT_15,INIT_16,INIT_17,
		INIT_18,INIT_19,INIT_1A,INIT_1B,INIT_1C,INIT_1D,INIT_1E,INIT_1F,
		INIT_20,INIT_21,INIT_22,INIT_23,INIT_24,INIT_25,INIT_26,INIT_27,
		INIT_28,INIT_29,INIT_2A,INIT_2B,INIT_2C,INIT_2D,INIT_2E,INIT_2F,
		INIT_30,INIT_31,INIT_32,INIT_33,INIT_34,INIT_35,INIT_36,INIT_37,
		INIT_38,INIT_39,INIT_3A,INIT_3B,INIT_3C,INIT_3D,INIT_3E,INIT_3F : bit_vector
	);
	port(
		DO   : out std_logic_vector(15 downto 0);	-- Port 16-bit Data Output
		DOP  : out std_logic_vector(1  downto 0);	-- Port 2-bit Parity Output
		ADDR : in  std_logic_vector(9  downto 0); 	-- Port 10-bit Address Input
		CLK  : in  std_logic;			 			-- Port Clock
		DI   : in  std_logic_vector(15 downto 0); 	-- Port 16-bit Data Input
		DIP  : in  std_logic_vector(1  downto 0); 	-- Port 2-bit parity Input
		EN   : in  std_logic;			 			-- Port RAM Enable Input
		SSR  : in  std_logic;			 			-- Port Synchronous Set/Reset Input
		WE   : in  std_logic			 			-- Port Write Enable Input
	);
	end component;

begin

	addrin <= addr;
	clkin  <= clk;
	dout   <= doutout;

	-- FRAME0002_RAMB06 instantiation
	FRAME0002_RAMB06 : RAMB16_S18
	generic map (

		-- The following generics are only necessary if you wish to change the default behavior.
		WRITE_MODE => "NO_CHANGE", 	-- WRITE_FIRST, READ_FIRST or NO_CHANGE

		-- The following generic INIT_xx declarations are only necessary
		-- if you wish to change the initial contents of the RAM to anything
		-- other than all zero's.
		INIT_00 => x"51A4ED7857F3C2C237378034B4C38028A3A627D459FDF8DA335FBC4A9D66215C",
		INIT_01 => x"27CC7F0612285DC18A45D12E45CCDD7CA8C6174B1B7B3022E18AAADC642EE5FE",
		INIT_02 => x"34366C8E9B427DBB5C023AD3D35D211AF24D130B033B30025A760C485E0B46D4",
		INIT_03 => x"A5EB53361AAE5AB0516036ED65F1C43734B317A2A882A00C51A1CB6ACCC4E64B",
		INIT_04 => x"0F4CE16B46350A21D9CA41D2C1F169B9604E964E5830982C2AF0DCF5242B924C",
		INIT_05 => x"DE8455CC5AD493F8AD4FA8B60E213E8EC0FDF903C60C91EA0AB1A5E8685A9468",
		INIT_06 => x"00C6468CD0A04E7BDE47A565CA4E75D1BD74F8CA79A55C4E203DAEEC89E52572",
		INIT_07 => x"77D6CB8007FA55E14C6C18D0703011E00C97511EC34A8AA01FF97AC467EC34A6",
		INIT_08 => x"EE7F5817DAAA2AAF5247A24440CD5C8EBAD1879A441B116296A6CAED25A2CAA3",
		INIT_09 => x"2B68CE5FB50D6349FD1D6087CE068A6FA02D4D37C23F32FE41895AFC4CFD1B46",
		INIT_0A => x"CF806E3427126D66BCD050A8BF49266454810657D326161211537B67BCC06BDB",
		INIT_0B => x"FD2A8DA47EAE47ADBAE8F2F8B3943B7F4AA0D9904E31CE4DD2C5D9B1913E9323",
		INIT_0C => x"8A14FF645DAB1188978275171721060927D63720FB5E54B41F7134F8DA254CF5",
		INIT_0D => x"1056C967C5625CF119219D51671D0FF8D86BD46DB76AD6171800D59483FA42B7",
		INIT_0E => x"BD8565AE319C3510603974491E01332A91D5BA8C6D8E2050DC07359376092E87",
		INIT_0F => x"2D5B0D0B60B40554522270DA62F5859BAA694217B762AE1D97FA1D9939C64DCD",
		INIT_10 => x"32682794951541621CEA7F3D5C1E4F7C05023B8208C026E7EBBAA31762B197CD",
		INIT_11 => x"3E9F959685D233FFE76B3AA37938117187C7264872389A8199276BE5B84E6F9C",
		INIT_12 => x"E2A9C5669C61FD89057767A38FC5BDA7AB58ADC5C60EC36BECBC4A7A67BA3DEA",
		INIT_13 => x"0F70397CE90707BFE4185B54EB6132C0E65E8F56D392C5E76D43FBBEA75144A0",
		INIT_14 => x"79FEB6BB124C1BBD1588288B45EDF155CD80F3C24519095BA98481B77BFC4208",
		INIT_15 => x"783C689EEBAA24F82A745573C3FF197F50D7EF5FB681AA35675F49FE644E4982",
		INIT_16 => x"E77F49C1A00FCA05C1D6740CB319D698A966234CDD3413F6E76F29907F06B394",
		INIT_17 => x"22EF4A1D4069D6A140EABCFD781A3CCAA79B5A79DFD7AFAC60FDCC76904509B3",
		INIT_18 => x"4C82C27E8DAAB3D9F98F99BD206633397F954473C702F19868342EB58A432221",
		INIT_19 => x"0ADF485724FAE703FB123CB25821A11BC1546242F9A253A663BD7A55CF03B126",
		INIT_1A => x"375D78A4806DA34B0487BF1426E784F036142BD4BD1FDB260DE54266FD3148B4",
		INIT_1B => x"B0848F3443A9C67E56115848166B2D481504C27DE3F93F10B779823BA2DB389A",
		INIT_1C => x"3CD7E3CB7CB21D12915C7AFC9006D8D67CD7E23216CA0B024610D41C17ED62E0",
		INIT_1D => x"CD321567A94D6FCEE82ACD62DC53069AEBAB3929A0F3534D47D150CA7B501D18",
		INIT_1E => x"CBE431BB2D3A4862F41A4F1CA193D973272DFDF8C61720D50FDD0D48AC0714AA",
		INIT_1F => x"0DB0031EF3325EBB72BFB4EE5BBD92A36692BDA8253049EB292988827DFC0A55",
		INIT_20 => x"04F34F6AD4139923835DCD92CC620A166F0B88FC5B726F28A29E2B81AA191241",
		INIT_21 => x"DF51A77509A43A069B896F74C12E7F9F211DA692664D71F4548B454D7A988363",
		INIT_22 => x"3FDC79A799C29E937613C7CCAD3D0D0AB239BA0F558846D786A344E754F7EF39",
		INIT_23 => x"E7D7D9F2EF21717EE853C835F48E04B7F987FFF84112F943B18E83BD5ED2CC4F",
		INIT_24 => x"0F27C54C55D0C17EF5A38DAF07186AA28508A3596093D3E6527E06D401C8DBB1",
		INIT_25 => x"07DAD8252BE565436F98571AB620FFE8E365630E168DC84AB4483954C4E4E60B",
		INIT_26 => x"E44D3A6F1B021FF183B27662E7B249F11716C5BC11EEE5B5E118027AD6FC319A",
		INIT_27 => x"9E3F5ABA1A4D50BB33714411D0947871CA38B0D1F1BAC2FBAAFBD1548196A219",
		INIT_28 => x"3E78B307CB871C2C1E57CE22430C65CCB573A3329F6240B5DBEF0AF542BD4CDA",
		INIT_29 => x"2DBB834E24AD3C929D3760557998095C41EF5CC80ED9F9CB3243A9C5F6068ED8",
		INIT_2A => x"FB783245601CE6ACEF58E3C30C448FB7B88EE7A6407BB017E3AF4A255DA24630",
		INIT_2B => x"026C51BFCB368FA3F406A4C1819C5CB21C521C46E8694375ABCDD2B4A0325AB2",
		INIT_2C => x"73674DBD26DF3E868C1DA3C5C96CF8B7E85D90950C4E109A11E8503FE03FB051",
		INIT_2D => x"B8DA86005ACD1C4DEBA647B7B6D814B1EDA992A8C42EC29E966964734FDAA23A",
		INIT_2E => x"42AEE583E8C3B47BA642D6CFCDFF00F63FD3DB6DF4C30A15502EDB514DB9C8EB",
		INIT_2F => x"F3B8F3AB9BF89D046686B10655EA1EE88F3423F50ADB49DC4FC5CB495C3FDACF",
		INIT_30 => x"92DF22191F741A37F42EA4DE498FB4E856E6195A91303A2F4627BF7217C789C7",
		INIT_31 => x"5E7EE79FD592E753A6F9DBFE67B4A5A283447C44DFB7E1D82A49EA07CEB655D1",
		INIT_32 => x"3DEE703434B279436B683A492213CD543D433333F3DD283C4CB792C551086612",
		INIT_33 => x"53D63279A55EC478AD380DFFD998B65BE1054177DBB41B0261197F1CECE043D0",
		INIT_34 => x"FB55CB37C0E1353ED20BA4581701AFEB461C144AB8F9346A3F56EBC3ED9F15E7",
		INIT_35 => x"201E4E3F73AEC94BCECC0EEB546D6732542BE0C7EB9612F837A869B9974DFDE8",
		INIT_36 => x"C3DE992AEFF92EF4D95CE6B4502B7C5C9D12F4BBF8496C413DBF93C443813F55",
		INIT_37 => x"6048C88472C469153017D9DED7C7C40B4D54A6FBDB3527B30A1D824DB3DC6BC7",
		INIT_38 => x"626C668333C9D5DE9DC3DF5D05695E53170D6641E229760897B198AA9ED400D9",
		INIT_39 => x"92698FAE7B3D69F472F2410C00808366B391CD3D3287EFAECE24D98983A46917",
		INIT_3A => x"F7B009565AF77313970F1A1E3F3439BF8EA85E835A42CC53CD83058EEFCC80B9",
		INIT_3B => x"C43200DE2F088B49470D860E6000463FAAC40B55FEBB16FD8C91295A91988E53",
		INIT_3C => x"72C86F84A80EDD5E186EBAFF01A4A2C01CC5CE335A4A2D3FCBB1C1F82302A75D",
		INIT_3D => x"6FDF79366498C82EFD52DC1CECC1B0E3E214EDE0617BB101DF3F310253D8489F",
		INIT_3E => x"4FD50B459DD43F50DE797929091A2A16FA7324F185D2D154100E79ABE91999F7",
		INIT_3F => x"11111111111111111111111111111111C93B19B353900B8CA7492CCAD9FC4CD1"
	)port map (
		DO   => doutout,			-- Port 16-bit Data Output
		DOP  => open,				-- Port 2-bit Parity Output
		ADDR => addrin,				-- Port 10-bit Address Input
		CLK  => clkin, 				-- Port Clock
		DI   => (others => '0'),	-- Port 16-bit Data Input
		DIP  => (others => '0'),	-- Port 2-bit parity Input
		EN   => '1',				-- Port RAM Enable Input
		SSR  => '0',				-- Port Synchronous Set/Reset Input
		WE   => '0'					-- Port Write Enable Input
	);
	-- End of FRAME0002_RAMB06 instantiation

end FRAME0002_B2;